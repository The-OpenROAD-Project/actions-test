magic
tech sky130A
magscale 1 2
timestamp 1648858418
<< checkpaint >>
rect -3932 -3932 24449 26593
<< viali >>
rect 1409 19873 1443 19907
rect 2697 19873 2731 19907
rect 3157 19873 3191 19907
rect 6561 19873 6595 19907
rect 8953 19873 8987 19907
rect 11529 19873 11563 19907
rect 16681 19873 16715 19907
rect 18061 19873 18095 19907
rect 1685 19805 1719 19839
rect 3065 19805 3099 19839
rect 5457 19805 5491 19839
rect 6837 19805 6871 19839
rect 8033 19805 8067 19839
rect 9229 19805 9263 19839
rect 10425 19805 10459 19839
rect 10517 19805 10551 19839
rect 10609 19805 10643 19839
rect 10701 19805 10735 19839
rect 11805 19805 11839 19839
rect 13369 19805 13403 19839
rect 15853 19805 15887 19839
rect 16129 19805 16163 19839
rect 16957 19805 16991 19839
rect 18153 19805 18187 19839
rect 4353 19737 4387 19771
rect 7849 19737 7883 19771
rect 13553 19737 13587 19771
rect 14565 19737 14599 19771
rect 14749 19737 14783 19771
rect 4261 19669 4295 19703
rect 5365 19669 5399 19703
rect 10241 19669 10275 19703
rect 18521 19669 18555 19703
rect 8401 19465 8435 19499
rect 10977 19465 11011 19499
rect 11713 19465 11747 19499
rect 5365 19397 5399 19431
rect 9873 19397 9907 19431
rect 18429 19397 18463 19431
rect 1685 19329 1719 19363
rect 2973 19329 3007 19363
rect 4445 19329 4479 19363
rect 5273 19329 5307 19363
rect 5457 19329 5491 19363
rect 6745 19329 6779 19363
rect 7389 19329 7423 19363
rect 10149 19329 10183 19363
rect 10793 19329 10827 19363
rect 13461 19329 13495 19363
rect 13921 19329 13955 19363
rect 18705 19329 18739 19363
rect 1409 19261 1443 19295
rect 2697 19261 2731 19295
rect 4537 19261 4571 19295
rect 6561 19261 6595 19295
rect 6653 19261 6687 19295
rect 6837 19261 6871 19295
rect 10609 19261 10643 19295
rect 13185 19261 13219 19295
rect 14197 19261 14231 19295
rect 4721 19125 4755 19159
rect 6377 19125 6411 19159
rect 7481 19125 7515 19159
rect 15669 19125 15703 19159
rect 16957 19125 16991 19159
rect 1409 18921 1443 18955
rect 8033 18921 8067 18955
rect 10241 18921 10275 18955
rect 12449 18853 12483 18887
rect 3157 18785 3191 18819
rect 5825 18785 5859 18819
rect 6101 18785 6135 18819
rect 7573 18785 7607 18819
rect 8401 18785 8435 18819
rect 10701 18785 10735 18819
rect 12173 18785 12207 18819
rect 14657 18785 14691 18819
rect 14933 18785 14967 18819
rect 16037 18785 16071 18819
rect 16497 18785 16531 18819
rect 17785 18785 17819 18819
rect 3985 18717 4019 18751
rect 4077 18717 4111 18751
rect 4629 18717 4663 18751
rect 4813 18717 4847 18751
rect 8217 18717 8251 18751
rect 8953 18717 8987 18751
rect 9229 18717 9263 18751
rect 10609 18717 10643 18751
rect 11253 18717 11287 18751
rect 12081 18717 12115 18751
rect 12909 18717 12943 18751
rect 13093 18717 13127 18751
rect 15025 18717 15059 18751
rect 15853 18717 15887 18751
rect 16773 18717 16807 18751
rect 18061 18717 18095 18751
rect 2881 18649 2915 18683
rect 13001 18649 13035 18683
rect 3801 18581 3835 18615
rect 4629 18581 4663 18615
rect 11437 18581 11471 18615
rect 15669 18581 15703 18615
rect 2697 18377 2731 18411
rect 4077 18377 4111 18411
rect 6561 18377 6595 18411
rect 8953 18377 8987 18411
rect 12909 18377 12943 18411
rect 14381 18377 14415 18411
rect 5549 18309 5583 18343
rect 9597 18309 9631 18343
rect 13829 18309 13863 18343
rect 16037 18309 16071 18343
rect 2881 18241 2915 18275
rect 3157 18241 3191 18275
rect 5825 18241 5859 18275
rect 6377 18241 6411 18275
rect 7389 18241 7423 18275
rect 9045 18241 9079 18275
rect 9505 18241 9539 18275
rect 9689 18241 9723 18275
rect 10333 18241 10367 18275
rect 11713 18241 11747 18275
rect 12357 18241 12391 18275
rect 13001 18241 13035 18275
rect 13737 18241 13771 18275
rect 14657 18241 14691 18275
rect 14841 18241 14875 18275
rect 16681 18241 16715 18275
rect 2973 18173 3007 18207
rect 3065 18173 3099 18207
rect 7021 18173 7055 18207
rect 7481 18173 7515 18207
rect 10425 18173 10459 18207
rect 14565 18173 14599 18207
rect 14749 18173 14783 18207
rect 16957 18173 16991 18207
rect 12173 18105 12207 18139
rect 15853 18105 15887 18139
rect 10609 18037 10643 18071
rect 11529 18037 11563 18071
rect 18429 18037 18463 18071
rect 2145 17833 2179 17867
rect 5641 17833 5675 17867
rect 15301 17833 15335 17867
rect 17049 17833 17083 17867
rect 15945 17765 15979 17799
rect 2789 17697 2823 17731
rect 10701 17697 10735 17731
rect 12265 17697 12299 17731
rect 16773 17697 16807 17731
rect 16865 17697 16899 17731
rect 18705 17697 18739 17731
rect 2237 17629 2271 17663
rect 2881 17629 2915 17663
rect 4537 17629 4571 17663
rect 5181 17629 5215 17663
rect 5825 17629 5859 17663
rect 6285 17629 6319 17663
rect 6929 17629 6963 17663
rect 11345 17629 11379 17663
rect 12173 17629 12207 17663
rect 12357 17629 12391 17663
rect 12449 17629 12483 17663
rect 13001 17629 13035 17663
rect 13185 17629 13219 17663
rect 13369 17629 13403 17663
rect 14289 17629 14323 17663
rect 14473 17629 14507 17663
rect 15393 17629 15427 17663
rect 15853 17629 15887 17663
rect 16037 17629 16071 17663
rect 16589 17629 16623 17663
rect 16681 17629 16715 17663
rect 18429 17629 18463 17663
rect 10425 17561 10459 17595
rect 3249 17493 3283 17527
rect 4353 17493 4387 17527
rect 5089 17493 5123 17527
rect 6469 17493 6503 17527
rect 7113 17493 7147 17527
rect 8953 17493 8987 17527
rect 11161 17493 11195 17527
rect 11989 17493 12023 17527
rect 14381 17493 14415 17527
rect 8125 17289 8159 17323
rect 9229 17289 9263 17323
rect 13277 17289 13311 17323
rect 17141 17289 17175 17323
rect 3893 17221 3927 17255
rect 11805 17221 11839 17255
rect 2973 17153 3007 17187
rect 6377 17153 6411 17187
rect 9137 17153 9171 17187
rect 9965 17153 9999 17187
rect 11529 17153 11563 17187
rect 14473 17153 14507 17187
rect 15761 17153 15795 17187
rect 17325 17153 17359 17187
rect 17509 17153 17543 17187
rect 18337 17153 18371 17187
rect 3617 17085 3651 17119
rect 5365 17085 5399 17119
rect 6653 17085 6687 17119
rect 9781 17085 9815 17119
rect 14565 17085 14599 17119
rect 18245 17085 18279 17119
rect 17969 17017 18003 17051
rect 3157 16949 3191 16983
rect 10149 16949 10183 16983
rect 14749 16949 14783 16983
rect 15669 16949 15703 16983
rect 6009 16745 6043 16779
rect 12081 16745 12115 16779
rect 12541 16745 12575 16779
rect 14736 16745 14770 16779
rect 18705 16745 18739 16779
rect 3157 16609 3191 16643
rect 4077 16609 4111 16643
rect 5825 16609 5859 16643
rect 9689 16609 9723 16643
rect 9965 16609 9999 16643
rect 10609 16609 10643 16643
rect 10701 16609 10735 16643
rect 10885 16609 10919 16643
rect 13001 16609 13035 16643
rect 14473 16609 14507 16643
rect 16957 16609 16991 16643
rect 3985 16541 4019 16575
rect 4169 16541 4203 16575
rect 4261 16541 4295 16575
rect 5733 16541 5767 16575
rect 6837 16541 6871 16575
rect 6929 16541 6963 16575
rect 9597 16541 9631 16575
rect 10793 16541 10827 16575
rect 11897 16541 11931 16575
rect 12909 16541 12943 16575
rect 2881 16473 2915 16507
rect 17233 16473 17267 16507
rect 1409 16405 1443 16439
rect 3801 16405 3835 16439
rect 10425 16405 10459 16439
rect 16221 16405 16255 16439
rect 1869 16201 1903 16235
rect 3801 16201 3835 16235
rect 5641 16201 5675 16235
rect 9505 16201 9539 16235
rect 12725 16201 12759 16235
rect 14749 16201 14783 16235
rect 15393 16201 15427 16235
rect 17233 16201 17267 16235
rect 18061 16201 18095 16235
rect 8033 16133 8067 16167
rect 16037 16133 16071 16167
rect 1961 16065 1995 16099
rect 2605 16065 2639 16099
rect 3433 16065 3467 16099
rect 3617 16065 3651 16099
rect 4261 16065 4295 16099
rect 4445 16065 4479 16099
rect 5549 16065 5583 16099
rect 5733 16065 5767 16099
rect 6746 16065 6780 16099
rect 7757 16065 7791 16099
rect 10333 16065 10367 16099
rect 12817 16065 12851 16099
rect 13461 16065 13495 16099
rect 13921 16065 13955 16099
rect 14565 16065 14599 16099
rect 15209 16065 15243 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 17969 16065 18003 16099
rect 2697 15997 2731 16031
rect 2973 15997 3007 16031
rect 6561 15997 6595 16031
rect 6653 15997 6687 16031
rect 6837 15997 6871 16031
rect 10241 15997 10275 16031
rect 16773 15997 16807 16031
rect 9965 15929 9999 15963
rect 4353 15861 4387 15895
rect 6377 15861 6411 15895
rect 13369 15861 13403 15895
rect 14105 15861 14139 15895
rect 7389 15657 7423 15691
rect 9045 15657 9079 15691
rect 10333 15657 10367 15691
rect 13277 15657 13311 15691
rect 16957 15657 16991 15691
rect 2973 15521 3007 15555
rect 5457 15521 5491 15555
rect 7849 15521 7883 15555
rect 11529 15521 11563 15555
rect 14565 15521 14599 15555
rect 2881 15453 2915 15487
rect 5181 15453 5215 15487
rect 7757 15453 7791 15487
rect 9137 15453 9171 15487
rect 10241 15453 10275 15487
rect 10425 15453 10459 15487
rect 14473 15453 14507 15487
rect 15393 15453 15427 15487
rect 15577 15453 15611 15487
rect 16037 15453 16071 15487
rect 16865 15453 16899 15487
rect 17509 15453 17543 15487
rect 18337 15453 18371 15487
rect 18429 15453 18463 15487
rect 11805 15385 11839 15419
rect 18153 15385 18187 15419
rect 3249 15317 3283 15351
rect 6929 15317 6963 15351
rect 14105 15317 14139 15351
rect 15209 15317 15243 15351
rect 16221 15317 16255 15351
rect 17601 15317 17635 15351
rect 6929 15113 6963 15147
rect 12817 15113 12851 15147
rect 18429 15113 18463 15147
rect 11897 15045 11931 15079
rect 12081 15045 12115 15079
rect 13369 15045 13403 15079
rect 4629 14977 4663 15011
rect 5273 14977 5307 15011
rect 7113 14977 7147 15011
rect 7297 14977 7331 15011
rect 7757 14977 7791 15011
rect 10149 14977 10183 15011
rect 10333 14977 10367 15011
rect 12633 14977 12667 15011
rect 12817 14977 12851 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 15393 14977 15427 15011
rect 16681 14977 16715 15011
rect 8033 14909 8067 14943
rect 14197 14909 14231 14943
rect 14381 14909 14415 14943
rect 15485 14909 15519 14943
rect 16957 14909 16991 14943
rect 15025 14841 15059 14875
rect 4537 14773 4571 14807
rect 5181 14773 5215 14807
rect 9505 14773 9539 14807
rect 10241 14773 10275 14807
rect 13461 14773 13495 14807
rect 14013 14773 14047 14807
rect 6101 14569 6135 14603
rect 6929 14569 6963 14603
rect 7573 14569 7607 14603
rect 9045 14569 9079 14603
rect 14362 14569 14396 14603
rect 15853 14569 15887 14603
rect 16681 14569 16715 14603
rect 17969 14501 18003 14535
rect 2697 14433 2731 14467
rect 5549 14433 5583 14467
rect 10333 14433 10367 14467
rect 14105 14433 14139 14467
rect 16957 14433 16991 14467
rect 17141 14433 17175 14467
rect 18245 14433 18279 14467
rect 1869 14365 1903 14399
rect 2513 14365 2547 14399
rect 2605 14365 2639 14399
rect 2789 14365 2823 14399
rect 6285 14365 6319 14399
rect 6837 14365 6871 14399
rect 7481 14365 7515 14399
rect 9137 14365 9171 14399
rect 10425 14365 10459 14399
rect 11437 14365 11471 14399
rect 12357 14365 12391 14399
rect 13553 14365 13587 14399
rect 16865 14365 16899 14399
rect 17049 14365 17083 14399
rect 18337 14365 18371 14399
rect 1777 14297 1811 14331
rect 5273 14297 5307 14331
rect 2329 14229 2363 14263
rect 3801 14229 3835 14263
rect 10793 14229 10827 14263
rect 11529 14229 11563 14263
rect 12173 14229 12207 14263
rect 13369 14229 13403 14263
rect 4629 14025 4663 14059
rect 8125 14025 8159 14059
rect 15025 14025 15059 14059
rect 15853 14025 15887 14059
rect 16865 14025 16899 14059
rect 1685 13957 1719 13991
rect 3617 13957 3651 13991
rect 11805 13957 11839 13991
rect 13737 13957 13771 13991
rect 1409 13889 1443 13923
rect 3801 13889 3835 13923
rect 4813 13889 4847 13923
rect 6377 13889 6411 13923
rect 9413 13889 9447 13923
rect 10425 13889 10459 13923
rect 10517 13889 10551 13923
rect 10609 13889 10643 13923
rect 11529 13889 11563 13923
rect 13921 13889 13955 13923
rect 15117 13889 15151 13923
rect 15669 13889 15703 13923
rect 16681 13889 16715 13923
rect 3157 13821 3191 13855
rect 3985 13821 4019 13855
rect 9505 13821 9539 13855
rect 9781 13821 9815 13855
rect 10241 13821 10275 13855
rect 10701 13821 10735 13855
rect 6634 13685 6668 13719
rect 13277 13685 13311 13719
rect 2237 13481 2271 13515
rect 6101 13481 6135 13515
rect 6745 13481 6779 13515
rect 10057 13481 10091 13515
rect 14197 13481 14231 13515
rect 18705 13481 18739 13515
rect 7665 13413 7699 13447
rect 12541 13413 12575 13447
rect 2697 13345 2731 13379
rect 5917 13345 5951 13379
rect 11437 13345 11471 13379
rect 11529 13345 11563 13379
rect 16037 13345 16071 13379
rect 16957 13345 16991 13379
rect 2605 13277 2639 13311
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 5825 13277 5859 13311
rect 9689 13277 9723 13311
rect 9873 13277 9907 13311
rect 11345 13277 11379 13311
rect 11621 13277 11655 13311
rect 14105 13277 14139 13311
rect 14841 13277 14875 13311
rect 16129 13277 16163 13311
rect 6837 13209 6871 13243
rect 7849 13209 7883 13243
rect 12725 13209 12759 13243
rect 17233 13209 17267 13243
rect 3893 13141 3927 13175
rect 11161 13141 11195 13175
rect 14933 13141 14967 13175
rect 16497 13141 16531 13175
rect 4905 12937 4939 12971
rect 7481 12937 7515 12971
rect 8953 12937 8987 12971
rect 13369 12937 13403 12971
rect 15669 12937 15703 12971
rect 17785 12937 17819 12971
rect 18521 12937 18555 12971
rect 8309 12869 8343 12903
rect 9965 12869 9999 12903
rect 15577 12869 15611 12903
rect 2605 12801 2639 12835
rect 3985 12801 4019 12835
rect 4997 12801 5031 12835
rect 6561 12801 6595 12835
rect 6653 12801 6687 12835
rect 7389 12801 7423 12835
rect 7573 12801 7607 12835
rect 8125 12801 8159 12835
rect 8861 12801 8895 12835
rect 12725 12801 12759 12835
rect 13553 12801 13587 12835
rect 14749 12801 14783 12835
rect 17141 12801 17175 12835
rect 17325 12801 17359 12835
rect 17785 12801 17819 12835
rect 17969 12801 18003 12835
rect 18429 12801 18463 12835
rect 2513 12733 2547 12767
rect 6745 12733 6779 12767
rect 6837 12733 6871 12767
rect 9781 12733 9815 12767
rect 12357 12733 12391 12767
rect 12817 12733 12851 12767
rect 13737 12733 13771 12767
rect 2973 12665 3007 12699
rect 4077 12597 4111 12631
rect 6377 12597 6411 12631
rect 14933 12597 14967 12631
rect 6837 12393 6871 12427
rect 12633 12393 12667 12427
rect 3801 12257 3835 12291
rect 7297 12257 7331 12291
rect 11161 12257 11195 12291
rect 14565 12257 14599 12291
rect 16405 12257 16439 12291
rect 7205 12189 7239 12223
rect 10241 12189 10275 12223
rect 10425 12189 10459 12223
rect 10885 12189 10919 12223
rect 14841 12189 14875 12223
rect 16221 12189 16255 12223
rect 16313 12189 16347 12223
rect 16497 12189 16531 12223
rect 4077 12121 4111 12155
rect 7849 12121 7883 12155
rect 8033 12121 8067 12155
rect 5549 12053 5583 12087
rect 10333 12053 10367 12087
rect 16037 12053 16071 12087
rect 6929 11849 6963 11883
rect 8401 11849 8435 11883
rect 10701 11849 10735 11883
rect 11989 11849 12023 11883
rect 14473 11849 14507 11883
rect 4537 11781 4571 11815
rect 4721 11781 4755 11815
rect 9873 11781 9907 11815
rect 13553 11781 13587 11815
rect 1409 11713 1443 11747
rect 2513 11713 2547 11747
rect 5825 11713 5859 11747
rect 7113 11713 7147 11747
rect 10793 11713 10827 11747
rect 11897 11713 11931 11747
rect 12633 11713 12667 11747
rect 13369 11713 13403 11747
rect 13645 11713 13679 11747
rect 14289 11713 14323 11747
rect 14565 11713 14599 11747
rect 15025 11713 15059 11747
rect 16681 11713 16715 11747
rect 18061 11713 18095 11747
rect 7297 11645 7331 11679
rect 10149 11645 10183 11679
rect 17693 11645 17727 11679
rect 18153 11645 18187 11679
rect 12817 11577 12851 11611
rect 15209 11577 15243 11611
rect 1593 11509 1627 11543
rect 2421 11509 2455 11543
rect 5733 11509 5767 11543
rect 13645 11509 13679 11543
rect 14105 11509 14139 11543
rect 16773 11509 16807 11543
rect 1409 11305 1443 11339
rect 6561 11305 6595 11339
rect 17877 11305 17911 11339
rect 7573 11237 7607 11271
rect 5089 11169 5123 11203
rect 7113 11169 7147 11203
rect 10149 11169 10183 11203
rect 14105 11169 14139 11203
rect 15669 11169 15703 11203
rect 17417 11169 17451 11203
rect 18245 11169 18279 11203
rect 3157 11101 3191 11135
rect 4813 11101 4847 11135
rect 7205 11101 7239 11135
rect 8217 11101 8251 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 12357 11101 12391 11135
rect 13185 11101 13219 11135
rect 13277 11101 13311 11135
rect 14289 11101 14323 11135
rect 14473 11101 14507 11135
rect 18061 11101 18095 11135
rect 2881 11033 2915 11067
rect 11897 11033 11931 11067
rect 15945 11033 15979 11067
rect 8125 10965 8159 10999
rect 9321 10965 9355 10999
rect 12449 10965 12483 10999
rect 5825 10761 5859 10795
rect 6837 10761 6871 10795
rect 12725 10761 12759 10795
rect 16129 10761 16163 10795
rect 18705 10761 18739 10795
rect 8309 10693 8343 10727
rect 14197 10693 14231 10727
rect 15025 10693 15059 10727
rect 17233 10693 17267 10727
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 4721 10625 4755 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 9321 10625 9355 10659
rect 10609 10625 10643 10659
rect 11713 10625 11747 10659
rect 14933 10625 14967 10659
rect 15117 10625 15151 10659
rect 15761 10625 15795 10659
rect 4905 10557 4939 10591
rect 8585 10557 8619 10591
rect 9413 10557 9447 10591
rect 10517 10557 10551 10591
rect 11897 10557 11931 10591
rect 14473 10557 14507 10591
rect 15669 10557 15703 10591
rect 16957 10557 16991 10591
rect 9689 10489 9723 10523
rect 2973 10421 3007 10455
rect 4537 10421 4571 10455
rect 10885 10421 10919 10455
rect 11529 10421 11563 10455
rect 1869 10217 1903 10251
rect 5549 10217 5583 10251
rect 10701 10217 10735 10251
rect 11418 10217 11452 10251
rect 18061 10217 18095 10251
rect 1685 10081 1719 10115
rect 2973 10081 3007 10115
rect 6929 10081 6963 10115
rect 7113 10081 7147 10115
rect 8953 10081 8987 10115
rect 11161 10081 11195 10115
rect 15393 10081 15427 10115
rect 15485 10081 15519 10115
rect 1593 10013 1627 10047
rect 2881 10013 2915 10047
rect 3801 10013 3835 10047
rect 7021 10013 7055 10047
rect 7205 10013 7239 10047
rect 14749 10013 14783 10047
rect 15577 10013 15611 10047
rect 15669 10013 15703 10047
rect 17325 10013 17359 10047
rect 17969 10013 18003 10047
rect 4077 9945 4111 9979
rect 6193 9945 6227 9979
rect 9229 9945 9263 9979
rect 14565 9945 14599 9979
rect 3249 9877 3283 9911
rect 6101 9877 6135 9911
rect 6745 9877 6779 9911
rect 12909 9877 12943 9911
rect 15209 9877 15243 9911
rect 17417 9877 17451 9911
rect 1777 9673 1811 9707
rect 3893 9673 3927 9707
rect 9229 9673 9263 9707
rect 15669 9673 15703 9707
rect 6653 9605 6687 9639
rect 1685 9537 1719 9571
rect 1869 9537 1903 9571
rect 3617 9537 3651 9571
rect 4721 9537 4755 9571
rect 6377 9537 6411 9571
rect 9413 9537 9447 9571
rect 9505 9537 9539 9571
rect 10793 9537 10827 9571
rect 12817 9537 12851 9571
rect 15853 9537 15887 9571
rect 3433 9469 3467 9503
rect 3525 9469 3559 9503
rect 3709 9469 3743 9503
rect 4353 9469 4387 9503
rect 4813 9469 4847 9503
rect 9597 9469 9631 9503
rect 9689 9469 9723 9503
rect 10885 9469 10919 9503
rect 13461 9469 13495 9503
rect 13737 9469 13771 9503
rect 15209 9469 15243 9503
rect 16037 9469 16071 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 8125 9333 8159 9367
rect 10425 9333 10459 9367
rect 12633 9333 12667 9367
rect 18613 9333 18647 9367
rect 4169 9129 4203 9163
rect 7113 9129 7147 9163
rect 9965 9129 9999 9163
rect 13185 9129 13219 9163
rect 15485 9129 15519 9163
rect 16957 9129 16991 9163
rect 6561 9061 6595 9095
rect 7573 8993 7607 9027
rect 15209 8993 15243 9027
rect 17233 8993 17267 9027
rect 18521 8993 18555 9027
rect 4077 8925 4111 8959
rect 5641 8925 5675 8959
rect 6469 8925 6503 8959
rect 7481 8925 7515 8959
rect 10057 8925 10091 8959
rect 12081 8925 12115 8959
rect 14197 8925 14231 8959
rect 15117 8925 15151 8959
rect 16129 8925 16163 8959
rect 17141 8925 17175 8959
rect 17325 8925 17359 8959
rect 17417 8925 17451 8959
rect 18153 8925 18187 8959
rect 18337 8925 18371 8959
rect 4721 8857 4755 8891
rect 4905 8857 4939 8891
rect 13277 8857 13311 8891
rect 5549 8789 5583 8823
rect 11897 8789 11931 8823
rect 14289 8789 14323 8823
rect 15945 8789 15979 8823
rect 6561 8585 6595 8619
rect 7389 8585 7423 8619
rect 16681 8585 16715 8619
rect 3985 8517 4019 8551
rect 13277 8517 13311 8551
rect 14197 8517 14231 8551
rect 14841 8517 14875 8551
rect 16037 8517 16071 8551
rect 2053 8449 2087 8483
rect 2237 8449 2271 8483
rect 3065 8449 3099 8483
rect 3157 8449 3191 8483
rect 6377 8449 6411 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 8217 8449 8251 8483
rect 8401 8449 8435 8483
rect 10793 8449 10827 8483
rect 15945 8449 15979 8483
rect 16129 8449 16163 8483
rect 17049 8449 17083 8483
rect 18337 8449 18371 8483
rect 2145 8381 2179 8415
rect 2329 8381 2363 8415
rect 2881 8381 2915 8415
rect 3709 8381 3743 8415
rect 11805 8381 11839 8415
rect 13553 8381 13587 8415
rect 17141 8381 17175 8415
rect 17969 8381 18003 8415
rect 18429 8381 18463 8415
rect 5457 8313 5491 8347
rect 10885 8313 10919 8347
rect 14013 8313 14047 8347
rect 15025 8313 15059 8347
rect 1869 8245 1903 8279
rect 8309 8245 8343 8279
rect 6745 8041 6779 8075
rect 10701 8041 10735 8075
rect 13461 8041 13495 8075
rect 15853 8041 15887 8075
rect 1685 7905 1719 7939
rect 7573 7905 7607 7939
rect 7665 7905 7699 7939
rect 8953 7905 8987 7939
rect 12633 7905 12667 7939
rect 12909 7905 12943 7939
rect 14105 7905 14139 7939
rect 14381 7905 14415 7939
rect 1409 7837 1443 7871
rect 4813 7837 4847 7871
rect 5917 7837 5951 7871
rect 6653 7837 6687 7871
rect 7481 7837 7515 7871
rect 7758 7837 7792 7871
rect 13369 7837 13403 7871
rect 18245 7837 18279 7871
rect 9229 7769 9263 7803
rect 3157 7701 3191 7735
rect 4997 7701 5031 7735
rect 6009 7701 6043 7735
rect 7297 7701 7331 7735
rect 11161 7701 11195 7735
rect 18153 7701 18187 7735
rect 3341 7497 3375 7531
rect 9137 7497 9171 7531
rect 9965 7497 9999 7531
rect 10701 7497 10735 7531
rect 14841 7497 14875 7531
rect 15485 7497 15519 7531
rect 18705 7497 18739 7531
rect 6653 7429 6687 7463
rect 2605 7361 2639 7395
rect 3433 7361 3467 7395
rect 8769 7361 8803 7395
rect 10057 7361 10091 7395
rect 10793 7361 10827 7395
rect 13001 7361 13035 7395
rect 13093 7361 13127 7395
rect 13829 7361 13863 7395
rect 14933 7361 14967 7395
rect 15577 7361 15611 7395
rect 2237 7293 2271 7327
rect 2697 7293 2731 7327
rect 6377 7293 6411 7327
rect 8677 7293 8711 7327
rect 16957 7293 16991 7327
rect 17233 7293 17267 7327
rect 8125 7157 8159 7191
rect 12817 7157 12851 7191
rect 14013 7157 14047 7191
rect 7389 6953 7423 6987
rect 9597 6953 9631 6987
rect 17233 6885 17267 6919
rect 3801 6817 3835 6851
rect 7849 6817 7883 6851
rect 12449 6817 12483 6851
rect 12725 6817 12759 6851
rect 15853 6817 15887 6851
rect 16037 6817 16071 6851
rect 16773 6817 16807 6851
rect 7757 6749 7791 6783
rect 9781 6749 9815 6783
rect 12817 6749 12851 6783
rect 14841 6749 14875 6783
rect 15946 6749 15980 6783
rect 16129 6749 16163 6783
rect 16865 6749 16899 6783
rect 17693 6749 17727 6783
rect 17877 6749 17911 6783
rect 4077 6681 4111 6715
rect 17785 6681 17819 6715
rect 5549 6613 5583 6647
rect 14933 6613 14967 6647
rect 15669 6613 15703 6647
rect 3893 6409 3927 6443
rect 6469 6409 6503 6443
rect 7665 6409 7699 6443
rect 13277 6409 13311 6443
rect 16681 6409 16715 6443
rect 14197 6341 14231 6375
rect 1685 6273 1719 6307
rect 1869 6273 1903 6307
rect 4169 6273 4203 6307
rect 4261 6273 4295 6307
rect 5273 6273 5307 6307
rect 6377 6273 6411 6307
rect 7849 6273 7883 6307
rect 8033 6273 8067 6307
rect 13921 6273 13955 6307
rect 16865 6273 16899 6307
rect 17509 6273 17543 6307
rect 17693 6273 17727 6307
rect 4077 6205 4111 6239
rect 4353 6205 4387 6239
rect 5365 6205 5399 6239
rect 11529 6205 11563 6239
rect 11805 6205 11839 6239
rect 15669 6205 15703 6239
rect 17049 6205 17083 6239
rect 4905 6137 4939 6171
rect 1777 6069 1811 6103
rect 17601 6069 17635 6103
rect 3249 5865 3283 5899
rect 5089 5865 5123 5899
rect 8309 5865 8343 5899
rect 12357 5865 12391 5899
rect 15945 5865 15979 5899
rect 18705 5865 18739 5899
rect 5457 5729 5491 5763
rect 9505 5729 9539 5763
rect 12541 5729 12575 5763
rect 12817 5729 12851 5763
rect 15669 5729 15703 5763
rect 1501 5661 1535 5695
rect 4077 5661 4111 5695
rect 4261 5661 4295 5695
rect 5273 5661 5307 5695
rect 6561 5661 6595 5695
rect 9413 5661 9447 5695
rect 9597 5661 9631 5695
rect 9689 5661 9723 5695
rect 10701 5661 10735 5695
rect 10885 5661 10919 5695
rect 11069 5661 11103 5695
rect 12633 5661 12667 5695
rect 12725 5661 12759 5695
rect 15577 5661 15611 5695
rect 16957 5661 16991 5695
rect 1777 5593 1811 5627
rect 6837 5593 6871 5627
rect 17233 5593 17267 5627
rect 4169 5525 4203 5559
rect 9229 5525 9263 5559
rect 1501 5321 1535 5355
rect 3525 5321 3559 5355
rect 10885 5321 10919 5355
rect 17049 5321 17083 5355
rect 18337 5321 18371 5355
rect 9413 5253 9447 5287
rect 11621 5253 11655 5287
rect 13277 5253 13311 5287
rect 1869 5185 1903 5219
rect 3617 5185 3651 5219
rect 4261 5185 4295 5219
rect 6929 5185 6963 5219
rect 7113 5185 7147 5219
rect 8309 5185 8343 5219
rect 9137 5185 9171 5219
rect 11529 5185 11563 5219
rect 12357 5185 12391 5219
rect 13185 5185 13219 5219
rect 13369 5185 13403 5219
rect 14933 5185 14967 5219
rect 17417 5185 17451 5219
rect 18245 5185 18279 5219
rect 1961 5117 1995 5151
rect 4353 5117 4387 5151
rect 8401 5117 8435 5151
rect 12265 5117 12299 5151
rect 14749 5117 14783 5151
rect 17325 5117 17359 5151
rect 4629 5049 4663 5083
rect 12725 5049 12759 5083
rect 7021 4981 7055 5015
rect 8585 4981 8619 5015
rect 15117 4981 15151 5015
rect 7665 4777 7699 4811
rect 8309 4777 8343 4811
rect 10425 4777 10459 4811
rect 12633 4777 12667 4811
rect 6929 4709 6963 4743
rect 2237 4641 2271 4675
rect 2329 4641 2363 4675
rect 6653 4641 6687 4675
rect 10885 4641 10919 4675
rect 15025 4641 15059 4675
rect 17417 4641 17451 4675
rect 2145 4573 2179 4607
rect 2421 4573 2455 4607
rect 5273 4573 5307 4607
rect 6561 4573 6595 4607
rect 7573 4573 7607 4607
rect 8217 4573 8251 4607
rect 8401 4573 8435 4607
rect 10793 4573 10827 4607
rect 12541 4573 12575 4607
rect 13369 4573 13403 4607
rect 14289 4573 14323 4607
rect 14473 4573 14507 4607
rect 15117 4573 15151 4607
rect 17325 4573 17359 4607
rect 17509 4573 17543 4607
rect 17601 4573 17635 4607
rect 18153 4573 18187 4607
rect 9505 4505 9539 4539
rect 14381 4505 14415 4539
rect 1961 4437 1995 4471
rect 5181 4437 5215 4471
rect 9413 4437 9447 4471
rect 13461 4437 13495 4471
rect 15485 4437 15519 4471
rect 17141 4437 17175 4471
rect 18245 4437 18279 4471
rect 2237 4233 2271 4267
rect 14289 4233 14323 4267
rect 12817 4165 12851 4199
rect 16957 4165 16991 4199
rect 1961 4097 1995 4131
rect 2053 4097 2087 4131
rect 3065 4097 3099 4131
rect 5825 4097 5859 4131
rect 7481 4097 7515 4131
rect 8125 4097 8159 4131
rect 12541 4097 12575 4131
rect 15025 4097 15059 4131
rect 15301 4097 15335 4131
rect 3157 4029 3191 4063
rect 4077 4029 4111 4063
rect 5549 4029 5583 4063
rect 8309 4029 8343 4063
rect 15117 4029 15151 4063
rect 15209 4029 15243 4063
rect 16681 4029 16715 4063
rect 2697 3961 2731 3995
rect 7389 3893 7423 3927
rect 7941 3893 7975 3927
rect 14841 3893 14875 3927
rect 18429 3893 18463 3927
rect 3157 3689 3191 3723
rect 13001 3689 13035 3723
rect 14933 3689 14967 3723
rect 17693 3689 17727 3723
rect 7665 3621 7699 3655
rect 17233 3621 17267 3655
rect 1409 3553 1443 3587
rect 1685 3553 1719 3587
rect 6837 3553 6871 3587
rect 6929 3553 6963 3587
rect 7113 3553 7147 3587
rect 8125 3553 8159 3587
rect 8953 3553 8987 3587
rect 10425 3553 10459 3587
rect 10701 3553 10735 3587
rect 14657 3553 14691 3587
rect 15485 3553 15519 3587
rect 17969 3553 18003 3587
rect 7021 3485 7055 3519
rect 8033 3485 8067 3519
rect 14565 3485 14599 3519
rect 18061 3485 18095 3519
rect 12725 3417 12759 3451
rect 15761 3417 15795 3451
rect 6653 3349 6687 3383
rect 2605 3145 2639 3179
rect 8309 3145 8343 3179
rect 9781 3145 9815 3179
rect 14749 3145 14783 3179
rect 15945 3145 15979 3179
rect 17601 3145 17635 3179
rect 6837 3077 6871 3111
rect 13277 3077 13311 3111
rect 2697 3009 2731 3043
rect 6561 3009 6595 3043
rect 9873 3009 9907 3043
rect 12357 3009 12391 3043
rect 13001 3009 13035 3043
rect 15853 3009 15887 3043
rect 17785 3009 17819 3043
rect 17969 3009 18003 3043
rect 12541 2873 12575 2907
rect 14197 2601 14231 2635
rect 10609 2533 10643 2567
rect 14289 2397 14323 2431
rect 10425 2329 10459 2363
<< metal1 >>
rect 1104 20154 19412 20176
rect 1104 20102 4001 20154
rect 4053 20102 4065 20154
rect 4117 20102 4129 20154
rect 4181 20102 4193 20154
rect 4245 20102 4257 20154
rect 4309 20102 10104 20154
rect 10156 20102 10168 20154
rect 10220 20102 10232 20154
rect 10284 20102 10296 20154
rect 10348 20102 10360 20154
rect 10412 20102 16206 20154
rect 16258 20102 16270 20154
rect 16322 20102 16334 20154
rect 16386 20102 16398 20154
rect 16450 20102 16462 20154
rect 16514 20102 19412 20154
rect 1104 20080 19412 20102
rect 20162 19972 20168 19984
rect 13372 19944 20168 19972
rect 290 19864 296 19916
rect 348 19904 354 19916
rect 1397 19907 1455 19913
rect 1397 19904 1409 19907
rect 348 19876 1409 19904
rect 348 19864 354 19876
rect 1397 19873 1409 19876
rect 1443 19873 1455 19907
rect 1397 19867 1455 19873
rect 2685 19907 2743 19913
rect 2685 19873 2697 19907
rect 2731 19904 2743 19907
rect 2774 19904 2780 19916
rect 2731 19876 2780 19904
rect 2731 19873 2743 19876
rect 2685 19867 2743 19873
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 3878 19904 3884 19916
rect 3191 19876 3884 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 3878 19864 3884 19876
rect 3936 19864 3942 19916
rect 6546 19904 6552 19916
rect 6507 19876 6552 19904
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 7098 19864 7104 19916
rect 7156 19904 7162 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 7156 19876 8953 19904
rect 7156 19864 7162 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 8941 19867 8999 19873
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 11517 19907 11575 19913
rect 11517 19904 11529 19907
rect 9364 19876 11529 19904
rect 9364 19864 9370 19876
rect 11517 19873 11529 19876
rect 11563 19873 11575 19907
rect 11517 19867 11575 19873
rect 1578 19796 1584 19848
rect 1636 19836 1642 19848
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1636 19808 1685 19836
rect 1636 19796 1642 19808
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 3050 19836 3056 19848
rect 3011 19808 3056 19836
rect 1673 19799 1731 19805
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 5442 19836 5448 19848
rect 5403 19808 5448 19836
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 6178 19796 6184 19848
rect 6236 19836 6242 19848
rect 6825 19839 6883 19845
rect 6825 19836 6837 19839
rect 6236 19808 6837 19836
rect 6236 19796 6242 19808
rect 6825 19805 6837 19808
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7800 19808 8033 19836
rect 7800 19796 7806 19808
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 8662 19796 8668 19848
rect 8720 19836 8726 19848
rect 9217 19839 9275 19845
rect 9217 19836 9229 19839
rect 8720 19808 9229 19836
rect 8720 19796 8726 19808
rect 9217 19805 9229 19808
rect 9263 19805 9275 19839
rect 10410 19836 10416 19848
rect 10371 19808 10416 19836
rect 9217 19799 9275 19805
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19836 10747 19839
rect 10962 19836 10968 19848
rect 10735 19808 10968 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 4154 19728 4160 19780
rect 4212 19768 4218 19780
rect 4341 19771 4399 19777
rect 4341 19768 4353 19771
rect 4212 19740 4353 19768
rect 4212 19728 4218 19740
rect 4341 19737 4353 19740
rect 4387 19737 4399 19771
rect 4341 19731 4399 19737
rect 7558 19728 7564 19780
rect 7616 19768 7622 19780
rect 7837 19771 7895 19777
rect 7837 19768 7849 19771
rect 7616 19740 7849 19768
rect 7616 19728 7622 19740
rect 7837 19737 7849 19740
rect 7883 19737 7895 19771
rect 7837 19731 7895 19737
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10520 19768 10548 19799
rect 9916 19740 10548 19768
rect 10612 19768 10640 19799
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 13372 19845 13400 19944
rect 20162 19932 20168 19944
rect 20220 19932 20226 19984
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 15804 19876 16681 19904
rect 15804 19864 15810 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 17678 19904 17684 19916
rect 16669 19867 16727 19873
rect 16868 19876 17684 19904
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11756 19808 11805 19836
rect 11756 19796 11762 19808
rect 11793 19805 11805 19808
rect 11839 19805 11851 19839
rect 11793 19799 11851 19805
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 15562 19796 15568 19848
rect 15620 19836 15626 19848
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 15620 19808 15853 19836
rect 15620 19796 15626 19808
rect 15841 19805 15853 19808
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19836 16175 19839
rect 16868 19836 16896 19876
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 18046 19904 18052 19916
rect 18007 19876 18052 19904
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 16163 19808 16896 19836
rect 16945 19839 17003 19845
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 16945 19805 16957 19839
rect 16991 19836 17003 19839
rect 17126 19836 17132 19848
rect 16991 19808 17132 19836
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 18138 19836 18144 19848
rect 18099 19808 18144 19836
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 11054 19768 11060 19780
rect 10612 19740 11060 19768
rect 9916 19728 9922 19740
rect 11054 19728 11060 19740
rect 11112 19728 11118 19780
rect 13541 19771 13599 19777
rect 13541 19737 13553 19771
rect 13587 19768 13599 19771
rect 13630 19768 13636 19780
rect 13587 19740 13636 19768
rect 13587 19737 13599 19740
rect 13541 19731 13599 19737
rect 13630 19728 13636 19740
rect 13688 19728 13694 19780
rect 13998 19728 14004 19780
rect 14056 19768 14062 19780
rect 14553 19771 14611 19777
rect 14553 19768 14565 19771
rect 14056 19740 14565 19768
rect 14056 19728 14062 19740
rect 14553 19737 14565 19740
rect 14599 19737 14611 19771
rect 14553 19731 14611 19737
rect 14737 19771 14795 19777
rect 14737 19737 14749 19771
rect 14783 19768 14795 19771
rect 18230 19768 18236 19780
rect 14783 19740 18236 19768
rect 14783 19737 14795 19740
rect 14737 19731 14795 19737
rect 18230 19728 18236 19740
rect 18288 19728 18294 19780
rect 4249 19703 4307 19709
rect 4249 19669 4261 19703
rect 4295 19700 4307 19703
rect 4890 19700 4896 19712
rect 4295 19672 4896 19700
rect 4295 19669 4307 19672
rect 4249 19663 4307 19669
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 5074 19660 5080 19712
rect 5132 19700 5138 19712
rect 5353 19703 5411 19709
rect 5353 19700 5365 19703
rect 5132 19672 5365 19700
rect 5132 19660 5138 19672
rect 5353 19669 5365 19672
rect 5399 19669 5411 19703
rect 10226 19700 10232 19712
rect 10187 19672 10232 19700
rect 5353 19663 5411 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 18506 19700 18512 19712
rect 18467 19672 18512 19700
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 1104 19610 19412 19632
rect 1104 19558 7052 19610
rect 7104 19558 7116 19610
rect 7168 19558 7180 19610
rect 7232 19558 7244 19610
rect 7296 19558 7308 19610
rect 7360 19558 13155 19610
rect 13207 19558 13219 19610
rect 13271 19558 13283 19610
rect 13335 19558 13347 19610
rect 13399 19558 13411 19610
rect 13463 19558 19412 19610
rect 1104 19536 19412 19558
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 5442 19496 5448 19508
rect 5224 19468 5448 19496
rect 5224 19456 5230 19468
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 8389 19499 8447 19505
rect 8389 19465 8401 19499
rect 8435 19496 8447 19499
rect 10594 19496 10600 19508
rect 8435 19468 10600 19496
rect 8435 19465 8447 19468
rect 8389 19459 8447 19465
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 10962 19496 10968 19508
rect 10923 19468 10968 19496
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11701 19499 11759 19505
rect 11701 19465 11713 19499
rect 11747 19465 11759 19499
rect 16666 19496 16672 19508
rect 11701 19459 11759 19465
rect 13924 19468 16672 19496
rect 5353 19431 5411 19437
rect 5353 19428 5365 19431
rect 4448 19400 5365 19428
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 2961 19363 3019 19369
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 3326 19360 3332 19372
rect 3007 19332 3332 19360
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 4448 19369 4476 19400
rect 5353 19397 5365 19400
rect 5399 19397 5411 19431
rect 5460 19428 5488 19456
rect 5460 19400 7420 19428
rect 5353 19391 5411 19397
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5261 19363 5319 19369
rect 5261 19360 5273 19363
rect 4764 19332 5273 19360
rect 4764 19320 4770 19332
rect 5261 19329 5273 19332
rect 5307 19329 5319 19363
rect 5261 19323 5319 19329
rect 5445 19363 5503 19369
rect 5445 19329 5457 19363
rect 5491 19360 5503 19363
rect 5491 19332 6684 19360
rect 5491 19329 5503 19332
rect 5445 19323 5503 19329
rect 6656 19304 6684 19332
rect 6730 19320 6736 19372
rect 6788 19360 6794 19372
rect 7392 19369 7420 19400
rect 8846 19388 8852 19440
rect 8904 19388 8910 19440
rect 9861 19431 9919 19437
rect 9861 19397 9873 19431
rect 9907 19428 9919 19431
rect 10226 19428 10232 19440
rect 9907 19400 10232 19428
rect 9907 19397 9919 19400
rect 9861 19391 9919 19397
rect 10226 19388 10232 19400
rect 10284 19388 10290 19440
rect 7377 19363 7435 19369
rect 6788 19332 6833 19360
rect 6788 19320 6794 19332
rect 7377 19329 7389 19363
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 10137 19363 10195 19369
rect 10137 19329 10149 19363
rect 10183 19360 10195 19363
rect 10686 19360 10692 19372
rect 10183 19332 10692 19360
rect 10183 19329 10195 19332
rect 10137 19323 10195 19329
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 11716 19360 11744 19459
rect 12894 19428 12900 19440
rect 12742 19400 12900 19428
rect 12894 19388 12900 19400
rect 12952 19388 12958 19440
rect 13924 19369 13952 19468
rect 16666 19456 16672 19468
rect 16724 19496 16730 19508
rect 16724 19468 18736 19496
rect 16724 19456 16730 19468
rect 15194 19388 15200 19440
rect 15252 19388 15258 19440
rect 17954 19388 17960 19440
rect 18012 19388 18018 19440
rect 18417 19431 18475 19437
rect 18417 19397 18429 19431
rect 18463 19428 18475 19431
rect 18506 19428 18512 19440
rect 18463 19400 18512 19428
rect 18463 19397 18475 19400
rect 18417 19391 18475 19397
rect 18506 19388 18512 19400
rect 18564 19388 18570 19440
rect 18708 19369 18736 19468
rect 10836 19332 11744 19360
rect 13449 19363 13507 19369
rect 10836 19320 10842 19332
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 13909 19363 13967 19369
rect 13909 19360 13921 19363
rect 13495 19332 13921 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 13909 19329 13921 19332
rect 13955 19329 13967 19363
rect 13909 19323 13967 19329
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 842 19252 848 19304
rect 900 19292 906 19304
rect 1397 19295 1455 19301
rect 1397 19292 1409 19295
rect 900 19264 1409 19292
rect 900 19252 906 19264
rect 1397 19261 1409 19264
rect 1443 19261 1455 19295
rect 1397 19255 1455 19261
rect 2130 19252 2136 19304
rect 2188 19292 2194 19304
rect 2685 19295 2743 19301
rect 2685 19292 2697 19295
rect 2188 19264 2697 19292
rect 2188 19252 2194 19264
rect 2685 19261 2697 19264
rect 2731 19261 2743 19295
rect 2685 19255 2743 19261
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 6546 19292 6552 19304
rect 4571 19264 6552 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6825 19295 6883 19301
rect 6696 19264 6789 19292
rect 6696 19252 6702 19264
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 8018 19292 8024 19304
rect 6871 19264 8024 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 10594 19292 10600 19304
rect 10555 19264 10600 19292
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 12492 19264 13185 19292
rect 12492 19252 12498 19264
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 14182 19292 14188 19304
rect 14143 19264 14188 19292
rect 13173 19255 13231 19261
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 1486 19184 1492 19236
rect 1544 19224 1550 19236
rect 4154 19224 4160 19236
rect 1544 19196 4160 19224
rect 1544 19184 1550 19196
rect 4154 19184 4160 19196
rect 4212 19184 4218 19236
rect 5810 19184 5816 19236
rect 5868 19224 5874 19236
rect 6914 19224 6920 19236
rect 5868 19196 6920 19224
rect 5868 19184 5874 19196
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 3602 19156 3608 19168
rect 2924 19128 3608 19156
rect 2924 19116 2930 19128
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 4709 19159 4767 19165
rect 4709 19125 4721 19159
rect 4755 19156 4767 19159
rect 5534 19156 5540 19168
rect 4755 19128 5540 19156
rect 4755 19125 4767 19128
rect 4709 19119 4767 19125
rect 5534 19116 5540 19128
rect 5592 19116 5598 19168
rect 6086 19116 6092 19168
rect 6144 19156 6150 19168
rect 6365 19159 6423 19165
rect 6365 19156 6377 19159
rect 6144 19128 6377 19156
rect 6144 19116 6150 19128
rect 6365 19125 6377 19128
rect 6411 19125 6423 19159
rect 7466 19156 7472 19168
rect 7427 19128 7472 19156
rect 6365 19119 6423 19125
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 15654 19156 15660 19168
rect 15615 19128 15660 19156
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 16945 19159 17003 19165
rect 16945 19156 16957 19159
rect 15896 19128 16957 19156
rect 15896 19116 15902 19128
rect 16945 19125 16957 19128
rect 16991 19125 17003 19159
rect 16945 19119 17003 19125
rect 1104 19066 19412 19088
rect 1104 19014 4001 19066
rect 4053 19014 4065 19066
rect 4117 19014 4129 19066
rect 4181 19014 4193 19066
rect 4245 19014 4257 19066
rect 4309 19014 10104 19066
rect 10156 19014 10168 19066
rect 10220 19014 10232 19066
rect 10284 19014 10296 19066
rect 10348 19014 10360 19066
rect 10412 19014 16206 19066
rect 16258 19014 16270 19066
rect 16322 19014 16334 19066
rect 16386 19014 16398 19066
rect 16450 19014 16462 19066
rect 16514 19014 19412 19066
rect 1104 18992 19412 19014
rect 1397 18955 1455 18961
rect 1397 18921 1409 18955
rect 1443 18952 1455 18955
rect 3050 18952 3056 18964
rect 1443 18924 3056 18952
rect 1443 18921 1455 18924
rect 1397 18915 1455 18921
rect 3050 18912 3056 18924
rect 3108 18952 3114 18964
rect 8018 18952 8024 18964
rect 3108 18924 4108 18952
rect 7979 18924 8024 18952
rect 3108 18912 3114 18924
rect 4080 18896 4108 18924
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 10229 18955 10287 18961
rect 10229 18921 10241 18955
rect 10275 18952 10287 18955
rect 10502 18952 10508 18964
rect 10275 18924 10508 18952
rect 10275 18921 10287 18924
rect 10229 18915 10287 18921
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 16022 18952 16028 18964
rect 14608 18924 16028 18952
rect 14608 18912 14614 18924
rect 16022 18912 16028 18924
rect 16080 18912 16086 18964
rect 4062 18844 4068 18896
rect 4120 18844 4126 18896
rect 12434 18844 12440 18896
rect 12492 18884 12498 18896
rect 15838 18884 15844 18896
rect 12492 18856 12537 18884
rect 14936 18856 15844 18884
rect 12492 18844 12498 18856
rect 3145 18819 3203 18825
rect 3145 18785 3157 18819
rect 3191 18816 3203 18819
rect 5810 18816 5816 18828
rect 3191 18788 5816 18816
rect 3191 18785 3203 18788
rect 3145 18779 3203 18785
rect 5810 18776 5816 18788
rect 5868 18776 5874 18828
rect 6086 18816 6092 18828
rect 6047 18788 6092 18816
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 7432 18788 7573 18816
rect 7432 18776 7438 18788
rect 7561 18785 7573 18788
rect 7607 18816 7619 18819
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 7607 18788 8401 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 8389 18785 8401 18788
rect 8435 18785 8447 18819
rect 8389 18779 8447 18785
rect 10689 18819 10747 18825
rect 10689 18785 10701 18819
rect 10735 18816 10747 18819
rect 10778 18816 10784 18828
rect 10735 18788 10784 18816
rect 10735 18785 10747 18788
rect 10689 18779 10747 18785
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 12158 18816 12164 18828
rect 12119 18788 12164 18816
rect 12158 18776 12164 18788
rect 12216 18776 12222 18828
rect 14550 18776 14556 18828
rect 14608 18816 14614 18828
rect 14936 18825 14964 18856
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 14645 18819 14703 18825
rect 14645 18816 14657 18819
rect 14608 18788 14657 18816
rect 14608 18776 14614 18788
rect 14645 18785 14657 18788
rect 14691 18785 14703 18819
rect 14645 18779 14703 18785
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18785 14979 18819
rect 15654 18816 15660 18828
rect 14921 18779 14979 18785
rect 15028 18788 15660 18816
rect 3786 18708 3792 18760
rect 3844 18708 3850 18760
rect 3878 18708 3884 18760
rect 3936 18748 3942 18760
rect 3973 18751 4031 18757
rect 3973 18748 3985 18751
rect 3936 18720 3985 18748
rect 3936 18708 3942 18720
rect 3973 18717 3985 18720
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 4062 18708 4068 18760
rect 4120 18748 4126 18760
rect 4120 18720 4165 18748
rect 4120 18708 4126 18720
rect 4430 18708 4436 18760
rect 4488 18748 4494 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 4488 18720 4629 18748
rect 4488 18708 4494 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 4798 18748 4804 18760
rect 4759 18720 4804 18748
rect 4617 18711 4675 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 8202 18748 8208 18760
rect 8163 18720 8208 18748
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8352 18720 8953 18748
rect 8352 18708 8358 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18748 9275 18751
rect 9398 18748 9404 18760
rect 9263 18720 9404 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 10594 18748 10600 18760
rect 10555 18720 10600 18748
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 11241 18751 11299 18757
rect 11241 18717 11253 18751
rect 11287 18717 11299 18751
rect 11241 18711 11299 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 2130 18640 2136 18692
rect 2188 18640 2194 18692
rect 2866 18680 2872 18692
rect 2827 18652 2872 18680
rect 2866 18640 2872 18652
rect 2924 18640 2930 18692
rect 3804 18680 3832 18708
rect 5718 18680 5724 18692
rect 3804 18652 5724 18680
rect 5718 18640 5724 18652
rect 5776 18640 5782 18692
rect 7466 18680 7472 18692
rect 7314 18652 7472 18680
rect 7466 18640 7472 18652
rect 7524 18640 7530 18692
rect 9582 18640 9588 18692
rect 9640 18680 9646 18692
rect 11256 18680 11284 18711
rect 9640 18652 11284 18680
rect 12084 18680 12112 18711
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 12897 18751 12955 18757
rect 12897 18748 12909 18751
rect 12308 18720 12909 18748
rect 12308 18708 12314 18720
rect 12897 18717 12909 18720
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 14274 18748 14280 18760
rect 13127 18720 14280 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 15028 18757 15056 18788
rect 15654 18776 15660 18788
rect 15712 18816 15718 18828
rect 16025 18819 16083 18825
rect 16025 18816 16037 18819
rect 15712 18788 16037 18816
rect 15712 18776 15718 18788
rect 16025 18785 16037 18788
rect 16071 18785 16083 18819
rect 16025 18779 16083 18785
rect 16114 18776 16120 18828
rect 16172 18816 16178 18828
rect 16485 18819 16543 18825
rect 16485 18816 16497 18819
rect 16172 18788 16497 18816
rect 16172 18776 16178 18788
rect 16485 18785 16497 18788
rect 16531 18785 16543 18819
rect 16485 18779 16543 18785
rect 17034 18776 17040 18828
rect 17092 18816 17098 18828
rect 17773 18819 17831 18825
rect 17773 18816 17785 18819
rect 17092 18788 17785 18816
rect 17092 18776 17098 18788
rect 17773 18785 17785 18788
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 15013 18751 15071 18757
rect 15013 18717 15025 18751
rect 15059 18717 15071 18751
rect 15838 18748 15844 18760
rect 15799 18720 15844 18748
rect 15013 18711 15071 18717
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18748 16819 18751
rect 17586 18748 17592 18760
rect 16807 18720 17592 18748
rect 16807 18717 16819 18720
rect 16761 18711 16819 18717
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18748 18107 18751
rect 18322 18748 18328 18760
rect 18095 18720 18328 18748
rect 18095 18717 18107 18720
rect 18049 18711 18107 18717
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 12989 18683 13047 18689
rect 12989 18680 13001 18683
rect 12084 18652 13001 18680
rect 9640 18640 9646 18652
rect 12989 18649 13001 18652
rect 13035 18649 13047 18683
rect 12989 18643 13047 18649
rect 3142 18572 3148 18624
rect 3200 18612 3206 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3200 18584 3801 18612
rect 3200 18572 3206 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 4338 18572 4344 18624
rect 4396 18612 4402 18624
rect 4617 18615 4675 18621
rect 4617 18612 4629 18615
rect 4396 18584 4629 18612
rect 4396 18572 4402 18584
rect 4617 18581 4629 18584
rect 4663 18581 4675 18615
rect 4617 18575 4675 18581
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 11388 18584 11437 18612
rect 11388 18572 11394 18584
rect 11425 18581 11437 18584
rect 11471 18581 11483 18615
rect 11425 18575 11483 18581
rect 14826 18572 14832 18624
rect 14884 18612 14890 18624
rect 15657 18615 15715 18621
rect 15657 18612 15669 18615
rect 14884 18584 15669 18612
rect 14884 18572 14890 18584
rect 15657 18581 15669 18584
rect 15703 18581 15715 18615
rect 15657 18575 15715 18581
rect 1104 18522 19412 18544
rect 1104 18470 7052 18522
rect 7104 18470 7116 18522
rect 7168 18470 7180 18522
rect 7232 18470 7244 18522
rect 7296 18470 7308 18522
rect 7360 18470 13155 18522
rect 13207 18470 13219 18522
rect 13271 18470 13283 18522
rect 13335 18470 13347 18522
rect 13399 18470 13411 18522
rect 13463 18470 19412 18522
rect 1104 18448 19412 18470
rect 2685 18411 2743 18417
rect 2685 18377 2697 18411
rect 2731 18408 2743 18411
rect 2866 18408 2872 18420
rect 2731 18380 2872 18408
rect 2731 18377 2743 18380
rect 2685 18371 2743 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3878 18368 3884 18420
rect 3936 18408 3942 18420
rect 4065 18411 4123 18417
rect 4065 18408 4077 18411
rect 3936 18380 4077 18408
rect 3936 18368 3942 18380
rect 4065 18377 4077 18380
rect 4111 18377 4123 18411
rect 4065 18371 4123 18377
rect 4614 18368 4620 18420
rect 4672 18408 4678 18420
rect 6549 18411 6607 18417
rect 4672 18380 6408 18408
rect 4672 18368 4678 18380
rect 5074 18300 5080 18352
rect 5132 18300 5138 18352
rect 5534 18340 5540 18352
rect 5495 18312 5540 18340
rect 5534 18300 5540 18312
rect 5592 18300 5598 18352
rect 2774 18232 2780 18284
rect 2832 18272 2838 18284
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2832 18244 2881 18272
rect 2832 18232 2838 18244
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 3142 18272 3148 18284
rect 3103 18244 3148 18272
rect 2869 18235 2927 18241
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 5810 18232 5816 18284
rect 5868 18272 5874 18284
rect 6380 18281 6408 18380
rect 6549 18377 6561 18411
rect 6595 18408 6607 18411
rect 6638 18408 6644 18420
rect 6595 18380 6644 18408
rect 6595 18377 6607 18380
rect 6549 18371 6607 18377
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 8846 18368 8852 18420
rect 8904 18408 8910 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 8904 18380 8953 18408
rect 8904 18368 8910 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 8941 18371 8999 18377
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 12894 18408 12900 18420
rect 10008 18380 11008 18408
rect 12855 18380 12900 18408
rect 10008 18368 10014 18380
rect 9585 18343 9643 18349
rect 9585 18309 9597 18343
rect 9631 18340 9643 18343
rect 9631 18312 10364 18340
rect 9631 18309 9643 18312
rect 9585 18303 9643 18309
rect 6365 18275 6423 18281
rect 5868 18244 5913 18272
rect 5868 18232 5874 18244
rect 6365 18241 6377 18275
rect 6411 18241 6423 18275
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 6365 18235 6423 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18272 9091 18275
rect 9122 18272 9128 18284
rect 9079 18244 9128 18272
rect 9079 18241 9091 18244
rect 9033 18235 9091 18241
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 9858 18272 9864 18284
rect 9723 18244 9864 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18173 3019 18207
rect 2961 18167 3019 18173
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18204 3111 18207
rect 3099 18176 5764 18204
rect 3099 18173 3111 18176
rect 3053 18167 3111 18173
rect 2976 18068 3004 18167
rect 3602 18096 3608 18148
rect 3660 18136 3666 18148
rect 4522 18136 4528 18148
rect 3660 18108 4528 18136
rect 3660 18096 3666 18108
rect 4522 18096 4528 18108
rect 4580 18096 4586 18148
rect 5736 18136 5764 18176
rect 6546 18164 6552 18216
rect 6604 18204 6610 18216
rect 7009 18207 7067 18213
rect 7009 18204 7021 18207
rect 6604 18176 7021 18204
rect 6604 18164 6610 18176
rect 7009 18173 7021 18176
rect 7055 18173 7067 18207
rect 7009 18167 7067 18173
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 8202 18204 8208 18216
rect 7515 18176 8208 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 9508 18204 9536 18235
rect 9858 18232 9864 18244
rect 9916 18272 9922 18284
rect 10336 18281 10364 18312
rect 10321 18275 10379 18281
rect 9916 18244 10272 18272
rect 9916 18232 9922 18244
rect 9950 18204 9956 18216
rect 9508 18176 9956 18204
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 6730 18136 6736 18148
rect 5736 18108 6736 18136
rect 6730 18096 6736 18108
rect 6788 18096 6794 18148
rect 10244 18136 10272 18244
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10980 18272 11008 18380
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 14369 18411 14427 18417
rect 14369 18408 14381 18411
rect 14240 18380 14381 18408
rect 14240 18368 14246 18380
rect 14369 18377 14381 18380
rect 14415 18377 14427 18411
rect 18874 18408 18880 18420
rect 14369 18371 14427 18377
rect 16040 18380 18880 18408
rect 11422 18300 11428 18352
rect 11480 18340 11486 18352
rect 13817 18343 13875 18349
rect 11480 18312 12388 18340
rect 11480 18300 11486 18312
rect 12360 18281 12388 18312
rect 13817 18309 13829 18343
rect 13863 18340 13875 18343
rect 15194 18340 15200 18352
rect 13863 18312 15200 18340
rect 13863 18309 13875 18312
rect 13817 18303 13875 18309
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 16040 18349 16068 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 16025 18343 16083 18349
rect 16025 18309 16037 18343
rect 16071 18309 16083 18343
rect 16025 18303 16083 18309
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 16632 18312 17434 18340
rect 16632 18300 16638 18312
rect 11701 18275 11759 18281
rect 11701 18272 11713 18275
rect 10980 18244 11713 18272
rect 10321 18235 10379 18241
rect 11701 18241 11713 18244
rect 11747 18241 11759 18275
rect 11701 18235 11759 18241
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12952 18244 13001 18272
rect 12952 18232 12958 18244
rect 12989 18241 13001 18244
rect 13035 18272 13047 18275
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13035 18244 13737 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 14642 18272 14648 18284
rect 14603 18244 14648 18272
rect 13725 18235 13783 18241
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 14826 18272 14832 18284
rect 14787 18244 14832 18272
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 16666 18272 16672 18284
rect 16627 18244 16672 18272
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 10502 18204 10508 18216
rect 10459 18176 10508 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10870 18164 10876 18216
rect 10928 18204 10934 18216
rect 11238 18204 11244 18216
rect 10928 18176 11244 18204
rect 10928 18164 10934 18176
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 13906 18164 13912 18216
rect 13964 18164 13970 18216
rect 14550 18204 14556 18216
rect 14511 18176 14556 18204
rect 14550 18164 14556 18176
rect 14608 18164 14614 18216
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18204 14795 18207
rect 16114 18204 16120 18216
rect 14783 18176 16120 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 16114 18164 16120 18176
rect 16172 18164 16178 18216
rect 16942 18204 16948 18216
rect 16903 18176 16948 18204
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 10244 18108 12173 18136
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 13924 18136 13952 18164
rect 15194 18136 15200 18148
rect 13924 18108 15200 18136
rect 12161 18099 12219 18105
rect 15194 18096 15200 18108
rect 15252 18096 15258 18148
rect 15838 18136 15844 18148
rect 15799 18108 15844 18136
rect 15838 18096 15844 18108
rect 15896 18096 15902 18148
rect 4798 18068 4804 18080
rect 2976 18040 4804 18068
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10560 18040 10609 18068
rect 10560 18028 10566 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 11204 18040 11529 18068
rect 11204 18028 11210 18040
rect 11517 18037 11529 18040
rect 11563 18037 11575 18071
rect 11517 18031 11575 18037
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13906 18068 13912 18080
rect 12768 18040 13912 18068
rect 12768 18028 12774 18040
rect 13906 18028 13912 18040
rect 13964 18028 13970 18080
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 17034 18068 17040 18080
rect 15344 18040 17040 18068
rect 15344 18028 15350 18040
rect 17034 18028 17040 18040
rect 17092 18028 17098 18080
rect 18414 18068 18420 18080
rect 18375 18040 18420 18068
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 1104 17978 19412 18000
rect 1104 17926 4001 17978
rect 4053 17926 4065 17978
rect 4117 17926 4129 17978
rect 4181 17926 4193 17978
rect 4245 17926 4257 17978
rect 4309 17926 10104 17978
rect 10156 17926 10168 17978
rect 10220 17926 10232 17978
rect 10284 17926 10296 17978
rect 10348 17926 10360 17978
rect 10412 17926 16206 17978
rect 16258 17926 16270 17978
rect 16322 17926 16334 17978
rect 16386 17926 16398 17978
rect 16450 17926 16462 17978
rect 16514 17926 19412 17978
rect 1104 17904 19412 17926
rect 2130 17864 2136 17876
rect 2091 17836 2136 17864
rect 2130 17824 2136 17836
rect 2188 17824 2194 17876
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 4856 17836 5641 17864
rect 4856 17824 4862 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 15289 17867 15347 17873
rect 15289 17833 15301 17867
rect 15335 17864 15347 17867
rect 16574 17864 16580 17876
rect 15335 17836 16580 17864
rect 15335 17833 15347 17836
rect 15289 17827 15347 17833
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 17037 17867 17095 17873
rect 17037 17864 17049 17867
rect 17000 17836 17049 17864
rect 17000 17824 17006 17836
rect 17037 17833 17049 17836
rect 17083 17833 17095 17867
rect 17037 17827 17095 17833
rect 15933 17799 15991 17805
rect 15933 17765 15945 17799
rect 15979 17796 15991 17799
rect 18230 17796 18236 17808
rect 15979 17768 18236 17796
rect 15979 17765 15991 17768
rect 15933 17759 15991 17765
rect 18230 17756 18236 17768
rect 18288 17756 18294 17808
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 10686 17728 10692 17740
rect 5592 17700 6316 17728
rect 10647 17700 10692 17728
rect 5592 17688 5598 17700
rect 1946 17620 1952 17672
rect 2004 17660 2010 17672
rect 2225 17663 2283 17669
rect 2225 17660 2237 17663
rect 2004 17632 2237 17660
rect 2004 17620 2010 17632
rect 2225 17629 2237 17632
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 2869 17663 2927 17669
rect 2869 17629 2881 17663
rect 2915 17660 2927 17663
rect 4338 17660 4344 17672
rect 2915 17632 4344 17660
rect 2915 17629 2927 17632
rect 2869 17623 2927 17629
rect 4338 17620 4344 17632
rect 4396 17620 4402 17672
rect 4522 17660 4528 17672
rect 4483 17632 4528 17660
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5718 17620 5724 17672
rect 5776 17660 5782 17672
rect 6288 17669 6316 17700
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 12250 17728 12256 17740
rect 12211 17700 12256 17728
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 15102 17728 15108 17740
rect 14292 17700 15108 17728
rect 14292 17672 14320 17700
rect 15102 17688 15108 17700
rect 15160 17728 15166 17740
rect 16761 17731 16819 17737
rect 16761 17728 16773 17731
rect 15160 17700 15884 17728
rect 15160 17688 15166 17700
rect 5813 17663 5871 17669
rect 5813 17660 5825 17663
rect 5776 17632 5825 17660
rect 5776 17620 5782 17632
rect 5813 17629 5825 17632
rect 5859 17629 5871 17663
rect 5813 17623 5871 17629
rect 6273 17663 6331 17669
rect 6273 17629 6285 17663
rect 6319 17629 6331 17663
rect 6914 17660 6920 17672
rect 6875 17632 6920 17660
rect 6273 17623 6331 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 9306 17620 9312 17672
rect 9364 17620 9370 17672
rect 11238 17620 11244 17672
rect 11296 17660 11302 17672
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 11296 17632 11345 17660
rect 11296 17620 11302 17632
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 12158 17660 12164 17672
rect 12119 17632 12164 17660
rect 11333 17623 11391 17629
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12989 17663 13047 17669
rect 12989 17660 13001 17663
rect 12483 17632 13001 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 12989 17629 13001 17632
rect 13035 17629 13047 17663
rect 12989 17623 13047 17629
rect 10413 17595 10471 17601
rect 10413 17561 10425 17595
rect 10459 17592 10471 17595
rect 10502 17592 10508 17604
rect 10459 17564 10508 17592
rect 10459 17561 10471 17564
rect 10413 17555 10471 17561
rect 10502 17552 10508 17564
rect 10560 17552 10566 17604
rect 10962 17552 10968 17604
rect 11020 17592 11026 17604
rect 12360 17592 12388 17623
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 13136 17632 13185 17660
rect 13136 17620 13142 17632
rect 13173 17629 13185 17632
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 13538 17660 13544 17672
rect 13403 17632 13544 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 14274 17660 14280 17672
rect 14235 17632 14280 17660
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14642 17660 14648 17672
rect 14507 17632 14648 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 14642 17620 14648 17632
rect 14700 17620 14706 17672
rect 15378 17660 15384 17672
rect 15339 17632 15384 17660
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 15856 17669 15884 17700
rect 16040 17700 16773 17728
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15930 17620 15936 17672
rect 15988 17660 15994 17672
rect 16040 17669 16068 17700
rect 16761 17697 16773 17700
rect 16807 17697 16819 17731
rect 16761 17691 16819 17697
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 18046 17728 18052 17740
rect 16899 17700 18052 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 18693 17731 18751 17737
rect 18693 17697 18705 17731
rect 18739 17728 18751 17731
rect 19518 17728 19524 17740
rect 18739 17700 19524 17728
rect 18739 17697 18751 17700
rect 18693 17691 18751 17697
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 16025 17663 16083 17669
rect 16025 17660 16037 17663
rect 15988 17632 16037 17660
rect 15988 17620 15994 17632
rect 16025 17629 16037 17632
rect 16071 17629 16083 17663
rect 16574 17660 16580 17672
rect 16535 17632 16580 17660
rect 16025 17623 16083 17629
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17629 16727 17663
rect 16669 17623 16727 17629
rect 11020 17564 12388 17592
rect 11020 17552 11026 17564
rect 16114 17552 16120 17604
rect 16172 17592 16178 17604
rect 16684 17592 16712 17623
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 18417 17663 18475 17669
rect 18417 17660 18429 17663
rect 18196 17632 18429 17660
rect 18196 17620 18202 17632
rect 18417 17629 18429 17632
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 17310 17592 17316 17604
rect 16172 17564 17316 17592
rect 16172 17552 16178 17564
rect 17310 17552 17316 17564
rect 17368 17552 17374 17604
rect 3237 17527 3295 17533
rect 3237 17493 3249 17527
rect 3283 17524 3295 17527
rect 3878 17524 3884 17536
rect 3283 17496 3884 17524
rect 3283 17493 3295 17496
rect 3237 17487 3295 17493
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4430 17524 4436 17536
rect 4387 17496 4436 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 5077 17527 5135 17533
rect 5077 17524 5089 17527
rect 5040 17496 5089 17524
rect 5040 17484 5046 17496
rect 5077 17493 5089 17496
rect 5123 17493 5135 17527
rect 5077 17487 5135 17493
rect 6457 17527 6515 17533
rect 6457 17493 6469 17527
rect 6503 17524 6515 17527
rect 6638 17524 6644 17536
rect 6503 17496 6644 17524
rect 6503 17493 6515 17496
rect 6457 17487 6515 17493
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 7101 17527 7159 17533
rect 7101 17493 7113 17527
rect 7147 17524 7159 17527
rect 7650 17524 7656 17536
rect 7147 17496 7656 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 8941 17527 8999 17533
rect 8941 17493 8953 17527
rect 8987 17524 8999 17527
rect 9674 17524 9680 17536
rect 8987 17496 9680 17524
rect 8987 17493 8999 17496
rect 8941 17487 8999 17493
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 10836 17496 11161 17524
rect 10836 17484 10842 17496
rect 11149 17493 11161 17496
rect 11195 17493 11207 17527
rect 11149 17487 11207 17493
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 11977 17527 12035 17533
rect 11977 17524 11989 17527
rect 11848 17496 11989 17524
rect 11848 17484 11854 17496
rect 11977 17493 11989 17496
rect 12023 17493 12035 17527
rect 11977 17487 12035 17493
rect 14369 17527 14427 17533
rect 14369 17493 14381 17527
rect 14415 17524 14427 17527
rect 14458 17524 14464 17536
rect 14415 17496 14464 17524
rect 14415 17493 14427 17496
rect 14369 17487 14427 17493
rect 14458 17484 14464 17496
rect 14516 17484 14522 17536
rect 1104 17434 19412 17456
rect 1104 17382 7052 17434
rect 7104 17382 7116 17434
rect 7168 17382 7180 17434
rect 7232 17382 7244 17434
rect 7296 17382 7308 17434
rect 7360 17382 13155 17434
rect 13207 17382 13219 17434
rect 13271 17382 13283 17434
rect 13335 17382 13347 17434
rect 13399 17382 13411 17434
rect 13463 17382 19412 17434
rect 1104 17360 19412 17382
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 8202 17320 8208 17332
rect 8159 17292 8208 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9306 17320 9312 17332
rect 9263 17292 9312 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 13265 17323 13323 17329
rect 13265 17289 13277 17323
rect 13311 17320 13323 17323
rect 13538 17320 13544 17332
rect 13311 17292 13544 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16632 17292 17141 17320
rect 16632 17280 16638 17292
rect 17129 17289 17141 17292
rect 17175 17289 17187 17323
rect 17129 17283 17187 17289
rect 3878 17252 3884 17264
rect 3839 17224 3884 17252
rect 3878 17212 3884 17224
rect 3936 17212 3942 17264
rect 6914 17212 6920 17264
rect 6972 17252 6978 17264
rect 11790 17252 11796 17264
rect 6972 17224 7130 17252
rect 11751 17224 11796 17252
rect 6972 17212 6978 17224
rect 11790 17212 11796 17224
rect 11848 17212 11854 17264
rect 12802 17212 12808 17264
rect 12860 17212 12866 17264
rect 2958 17184 2964 17196
rect 2919 17156 2964 17184
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 4982 17144 4988 17196
rect 5040 17144 5046 17196
rect 5810 17144 5816 17196
rect 5868 17184 5874 17196
rect 6362 17184 6368 17196
rect 5868 17156 6368 17184
rect 5868 17144 5874 17156
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 9122 17184 9128 17196
rect 9083 17156 9128 17184
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9732 17156 9965 17184
rect 9732 17144 9738 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 11514 17184 11520 17196
rect 10744 17156 11520 17184
rect 10744 17144 10750 17156
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 14458 17184 14464 17196
rect 14419 17156 14464 17184
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 15436 17156 15761 17184
rect 15436 17144 15442 17156
rect 15749 17153 15761 17156
rect 15795 17184 15807 17187
rect 16942 17184 16948 17196
rect 15795 17156 16948 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17184 17555 17187
rect 18325 17187 18383 17193
rect 18325 17184 18337 17187
rect 17543 17156 18337 17184
rect 17543 17153 17555 17156
rect 17497 17147 17555 17153
rect 18325 17153 18337 17156
rect 18371 17184 18383 17187
rect 18414 17184 18420 17196
rect 18371 17156 18420 17184
rect 18371 17153 18383 17156
rect 18325 17147 18383 17153
rect 3602 17116 3608 17128
rect 3563 17088 3608 17116
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 3878 17076 3884 17128
rect 3936 17116 3942 17128
rect 5353 17119 5411 17125
rect 5353 17116 5365 17119
rect 3936 17088 5365 17116
rect 3936 17076 3942 17088
rect 5353 17085 5365 17088
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 5994 17076 6000 17128
rect 6052 17116 6058 17128
rect 6641 17119 6699 17125
rect 6641 17116 6653 17119
rect 6052 17088 6653 17116
rect 6052 17076 6058 17088
rect 6641 17085 6653 17088
rect 6687 17085 6699 17119
rect 9766 17116 9772 17128
rect 9727 17088 9772 17116
rect 6641 17079 6699 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 14550 17116 14556 17128
rect 14511 17088 14556 17116
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 17328 17116 17356 17147
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 18230 17116 18236 17128
rect 17328 17088 18236 17116
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 17957 17051 18015 17057
rect 17957 17017 17969 17051
rect 18003 17048 18015 17051
rect 18046 17048 18052 17060
rect 18003 17020 18052 17048
rect 18003 17017 18015 17020
rect 17957 17011 18015 17017
rect 18046 17008 18052 17020
rect 18104 17008 18110 17060
rect 3145 16983 3203 16989
rect 3145 16949 3157 16983
rect 3191 16980 3203 16983
rect 4338 16980 4344 16992
rect 3191 16952 4344 16980
rect 3191 16949 3203 16952
rect 3145 16943 3203 16949
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 10137 16983 10195 16989
rect 10137 16949 10149 16983
rect 10183 16980 10195 16983
rect 10870 16980 10876 16992
rect 10183 16952 10876 16980
rect 10183 16949 10195 16952
rect 10137 16943 10195 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 14734 16980 14740 16992
rect 14695 16952 14740 16980
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 15746 16980 15752 16992
rect 15703 16952 15752 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 1104 16890 19412 16912
rect 1104 16838 4001 16890
rect 4053 16838 4065 16890
rect 4117 16838 4129 16890
rect 4181 16838 4193 16890
rect 4245 16838 4257 16890
rect 4309 16838 10104 16890
rect 10156 16838 10168 16890
rect 10220 16838 10232 16890
rect 10284 16838 10296 16890
rect 10348 16838 10360 16890
rect 10412 16838 16206 16890
rect 16258 16838 16270 16890
rect 16322 16838 16334 16890
rect 16386 16838 16398 16890
rect 16450 16838 16462 16890
rect 16514 16838 19412 16890
rect 1104 16816 19412 16838
rect 5994 16776 6000 16788
rect 5955 16748 6000 16776
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 12069 16779 12127 16785
rect 12069 16745 12081 16779
rect 12115 16776 12127 16779
rect 12250 16776 12256 16788
rect 12115 16748 12256 16776
rect 12115 16745 12127 16748
rect 12069 16739 12127 16745
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 14734 16785 14740 16788
rect 12529 16779 12587 16785
rect 12529 16776 12541 16779
rect 12406 16748 12541 16776
rect 5166 16668 5172 16720
rect 5224 16708 5230 16720
rect 10778 16708 10784 16720
rect 5224 16680 6868 16708
rect 5224 16668 5230 16680
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 3602 16640 3608 16652
rect 3191 16612 3608 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 3602 16600 3608 16612
rect 3660 16640 3666 16652
rect 3786 16640 3792 16652
rect 3660 16612 3792 16640
rect 3660 16600 3666 16612
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4338 16640 4344 16652
rect 4111 16612 4344 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 5813 16643 5871 16649
rect 4448 16612 5580 16640
rect 3970 16572 3976 16584
rect 3931 16544 3976 16572
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 1854 16464 1860 16516
rect 1912 16464 1918 16516
rect 2869 16507 2927 16513
rect 2869 16473 2881 16507
rect 2915 16473 2927 16507
rect 4172 16504 4200 16535
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 4304 16544 4349 16572
rect 4304 16532 4310 16544
rect 4448 16504 4476 16612
rect 5552 16516 5580 16612
rect 5813 16609 5825 16643
rect 5859 16640 5871 16643
rect 6546 16640 6552 16652
rect 5859 16612 6552 16640
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 5718 16572 5724 16584
rect 5679 16544 5724 16572
rect 5718 16532 5724 16544
rect 5776 16532 5782 16584
rect 6840 16581 6868 16680
rect 10704 16680 10784 16708
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10226 16640 10232 16652
rect 9999 16612 10232 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10226 16600 10232 16612
rect 10284 16640 10290 16652
rect 10704 16649 10732 16680
rect 10778 16668 10784 16680
rect 10836 16668 10842 16720
rect 12158 16668 12164 16720
rect 12216 16708 12222 16720
rect 12406 16708 12434 16748
rect 12529 16745 12541 16748
rect 12575 16745 12587 16779
rect 12529 16739 12587 16745
rect 14724 16779 14740 16785
rect 14724 16745 14736 16779
rect 14724 16739 14740 16745
rect 14734 16736 14740 16739
rect 14792 16736 14798 16788
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 18693 16779 18751 16785
rect 18693 16776 18705 16779
rect 18288 16748 18705 16776
rect 18288 16736 18294 16748
rect 18693 16745 18705 16748
rect 18739 16745 18751 16779
rect 18693 16739 18751 16745
rect 12216 16680 12434 16708
rect 12216 16668 12222 16680
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 10284 16612 10609 16640
rect 10284 16600 10290 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16609 10747 16643
rect 10870 16640 10876 16652
rect 10831 16612 10876 16640
rect 10689 16603 10747 16609
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 10962 16600 10968 16652
rect 11020 16600 11026 16652
rect 12986 16640 12992 16652
rect 12947 16612 12992 16640
rect 12986 16600 12992 16612
rect 13044 16600 13050 16652
rect 14461 16643 14519 16649
rect 14461 16609 14473 16643
rect 14507 16640 14519 16643
rect 16666 16640 16672 16652
rect 14507 16612 16672 16640
rect 14507 16609 14519 16612
rect 14461 16603 14519 16609
rect 16666 16600 16672 16612
rect 16724 16640 16730 16652
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16724 16612 16957 16640
rect 16724 16600 16730 16612
rect 16945 16609 16957 16612
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 6914 16532 6920 16584
rect 6972 16572 6978 16584
rect 9585 16575 9643 16581
rect 6972 16544 7017 16572
rect 6972 16532 6978 16544
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 9766 16572 9772 16584
rect 9631 16544 9772 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16572 10839 16575
rect 10980 16572 11008 16600
rect 10827 16544 11008 16572
rect 11885 16575 11943 16581
rect 10827 16541 10839 16544
rect 10781 16535 10839 16541
rect 11885 16541 11897 16575
rect 11931 16572 11943 16575
rect 12066 16572 12072 16584
rect 11931 16544 12072 16572
rect 11931 16541 11943 16544
rect 11885 16535 11943 16541
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 12897 16575 12955 16581
rect 12897 16541 12909 16575
rect 12943 16572 12955 16575
rect 13538 16572 13544 16584
rect 12943 16544 13544 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 5534 16504 5540 16516
rect 4172 16476 4476 16504
rect 5447 16476 5540 16504
rect 2869 16467 2927 16473
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 2590 16436 2596 16448
rect 1443 16408 2596 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 2590 16396 2596 16408
rect 2648 16396 2654 16448
rect 2884 16436 2912 16467
rect 5534 16464 5540 16476
rect 5592 16504 5598 16516
rect 6730 16504 6736 16516
rect 5592 16476 6736 16504
rect 5592 16464 5598 16476
rect 6730 16464 6736 16476
rect 6788 16464 6794 16516
rect 15746 16464 15752 16516
rect 15804 16464 15810 16516
rect 17218 16504 17224 16516
rect 17179 16476 17224 16504
rect 17218 16464 17224 16476
rect 17276 16464 17282 16516
rect 17678 16464 17684 16516
rect 17736 16464 17742 16516
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 2884 16408 3801 16436
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 8018 16396 8024 16448
rect 8076 16436 8082 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 8076 16408 10425 16436
rect 8076 16396 8082 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 16209 16439 16267 16445
rect 16209 16436 16221 16439
rect 15436 16408 16221 16436
rect 15436 16396 15442 16408
rect 16209 16405 16221 16408
rect 16255 16405 16267 16439
rect 16209 16399 16267 16405
rect 1104 16346 19412 16368
rect 1104 16294 7052 16346
rect 7104 16294 7116 16346
rect 7168 16294 7180 16346
rect 7232 16294 7244 16346
rect 7296 16294 7308 16346
rect 7360 16294 13155 16346
rect 13207 16294 13219 16346
rect 13271 16294 13283 16346
rect 13335 16294 13347 16346
rect 13399 16294 13411 16346
rect 13463 16294 19412 16346
rect 1104 16272 19412 16294
rect 1854 16232 1860 16244
rect 1815 16204 1860 16232
rect 1854 16192 1860 16204
rect 1912 16192 1918 16244
rect 3789 16235 3847 16241
rect 3789 16201 3801 16235
rect 3835 16232 3847 16235
rect 4246 16232 4252 16244
rect 3835 16204 4252 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 5718 16232 5724 16244
rect 5675 16204 5724 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5718 16192 5724 16204
rect 5776 16192 5782 16244
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 9493 16235 9551 16241
rect 6420 16204 6868 16232
rect 6420 16192 6426 16204
rect 6638 16164 6644 16176
rect 5736 16136 6644 16164
rect 1946 16096 1952 16108
rect 1907 16068 1952 16096
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 2590 16096 2596 16108
rect 2551 16068 2596 16096
rect 2590 16056 2596 16068
rect 2648 16096 2654 16108
rect 3421 16099 3479 16105
rect 3421 16096 3433 16099
rect 2648 16068 3433 16096
rect 2648 16056 2654 16068
rect 3421 16065 3433 16068
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 3878 16096 3884 16108
rect 3651 16068 3884 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 3878 16056 3884 16068
rect 3936 16056 3942 16108
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 4338 16096 4344 16108
rect 4295 16068 4344 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 4338 16056 4344 16068
rect 4396 16056 4402 16108
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 4614 16096 4620 16108
rect 4479 16068 4620 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 4614 16056 4620 16068
rect 4672 16096 4678 16108
rect 5736 16105 5764 16136
rect 6638 16124 6644 16136
rect 6696 16124 6702 16176
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 4672 16068 5549 16096
rect 4672 16056 4678 16068
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 5721 16099 5779 16105
rect 5721 16065 5733 16099
rect 5767 16065 5779 16099
rect 6730 16096 6736 16108
rect 6692 16068 6736 16096
rect 5721 16059 5779 16065
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 6840 16096 6868 16204
rect 9493 16201 9505 16235
rect 9539 16232 9551 16235
rect 9766 16232 9772 16244
rect 9539 16204 9772 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 12713 16235 12771 16241
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 12802 16232 12808 16244
rect 12759 16204 12808 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 14737 16235 14795 16241
rect 14737 16232 14749 16235
rect 14700 16204 14749 16232
rect 14700 16192 14706 16204
rect 14737 16201 14749 16204
rect 14783 16201 14795 16235
rect 14737 16195 14795 16201
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 15930 16232 15936 16244
rect 15427 16204 15936 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 17218 16232 17224 16244
rect 17179 16204 17224 16232
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 18012 16204 18061 16232
rect 18012 16192 18018 16204
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 8018 16164 8024 16176
rect 7979 16136 8024 16164
rect 8018 16124 8024 16136
rect 8076 16124 8082 16176
rect 9030 16124 9036 16176
rect 9088 16124 9094 16176
rect 13814 16124 13820 16176
rect 13872 16164 13878 16176
rect 13872 16136 14596 16164
rect 13872 16124 13878 16136
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 6840 16068 7757 16096
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 10502 16096 10508 16108
rect 10367 16068 10508 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16096 12863 16099
rect 12894 16096 12900 16108
rect 12851 16068 12900 16096
rect 12851 16065 12863 16068
rect 12805 16059 12863 16065
rect 12894 16056 12900 16068
rect 12952 16096 12958 16108
rect 13449 16099 13507 16105
rect 13449 16096 13461 16099
rect 12952 16068 13461 16096
rect 12952 16056 12958 16068
rect 13449 16065 13461 16068
rect 13495 16096 13507 16099
rect 13630 16096 13636 16108
rect 13495 16068 13636 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 13906 16096 13912 16108
rect 13867 16068 13912 16096
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 14568 16105 14596 16136
rect 15102 16124 15108 16176
rect 15160 16164 15166 16176
rect 16025 16167 16083 16173
rect 15160 16136 15976 16164
rect 15160 16124 15166 16136
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 15194 16096 15200 16108
rect 15155 16068 15200 16096
rect 14553 16059 14611 16065
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15948 16105 15976 16136
rect 16025 16133 16037 16167
rect 16071 16164 16083 16167
rect 16071 16136 16896 16164
rect 16071 16133 16083 16136
rect 16025 16127 16083 16133
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16574 16096 16580 16108
rect 16163 16068 16580 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 16868 16105 16896 16136
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 17494 16056 17500 16108
rect 17552 16096 17558 16108
rect 17957 16099 18015 16105
rect 17957 16096 17969 16099
rect 17552 16068 17969 16096
rect 17552 16056 17558 16068
rect 17957 16065 17969 16068
rect 18003 16065 18015 16099
rect 17957 16059 18015 16065
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 16028 2743 16031
rect 2958 16028 2964 16040
rect 2731 16000 2820 16028
rect 2871 16000 2964 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 2792 15960 2820 16000
rect 2958 15988 2964 16000
rect 3016 16028 3022 16040
rect 3970 16028 3976 16040
rect 3016 16000 3976 16028
rect 3016 15988 3022 16000
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 6546 16028 6552 16040
rect 6507 16000 6552 16028
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 6825 16031 6883 16037
rect 6696 16000 6741 16028
rect 6696 15988 6702 16000
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 6914 16028 6920 16040
rect 6871 16000 6920 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 10226 16028 10232 16040
rect 10187 16000 10232 16028
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 16761 16031 16819 16037
rect 16761 15997 16773 16031
rect 16807 16028 16819 16031
rect 16807 16000 16896 16028
rect 16807 15997 16819 16000
rect 16761 15991 16819 15997
rect 16868 15972 16896 16000
rect 3878 15960 3884 15972
rect 2792 15932 3884 15960
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 9214 15920 9220 15972
rect 9272 15960 9278 15972
rect 9953 15963 10011 15969
rect 9953 15960 9965 15963
rect 9272 15932 9965 15960
rect 9272 15920 9278 15932
rect 9953 15929 9965 15932
rect 9999 15929 10011 15963
rect 9953 15923 10011 15929
rect 16850 15920 16856 15972
rect 16908 15920 16914 15972
rect 4338 15892 4344 15904
rect 4299 15864 4344 15892
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 5442 15852 5448 15904
rect 5500 15892 5506 15904
rect 6365 15895 6423 15901
rect 6365 15892 6377 15895
rect 5500 15864 6377 15892
rect 5500 15852 5506 15864
rect 6365 15861 6377 15864
rect 6411 15861 6423 15895
rect 13354 15892 13360 15904
rect 13315 15864 13360 15892
rect 6365 15855 6423 15861
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14090 15892 14096 15904
rect 14051 15864 14096 15892
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 1104 15802 19412 15824
rect 1104 15750 4001 15802
rect 4053 15750 4065 15802
rect 4117 15750 4129 15802
rect 4181 15750 4193 15802
rect 4245 15750 4257 15802
rect 4309 15750 10104 15802
rect 10156 15750 10168 15802
rect 10220 15750 10232 15802
rect 10284 15750 10296 15802
rect 10348 15750 10360 15802
rect 10412 15750 16206 15802
rect 16258 15750 16270 15802
rect 16322 15750 16334 15802
rect 16386 15750 16398 15802
rect 16450 15750 16462 15802
rect 16514 15750 19412 15802
rect 1104 15728 19412 15750
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 7377 15691 7435 15697
rect 7377 15688 7389 15691
rect 6604 15660 7389 15688
rect 6604 15648 6610 15660
rect 7377 15657 7389 15660
rect 7423 15657 7435 15691
rect 9030 15688 9036 15700
rect 8991 15660 9036 15688
rect 7377 15651 7435 15657
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 10321 15691 10379 15697
rect 10321 15657 10333 15691
rect 10367 15688 10379 15691
rect 10502 15688 10508 15700
rect 10367 15660 10508 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 12986 15648 12992 15700
rect 13044 15688 13050 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 13044 15660 13277 15688
rect 13044 15648 13050 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 16945 15691 17003 15697
rect 16945 15657 16957 15691
rect 16991 15688 17003 15691
rect 17678 15688 17684 15700
rect 16991 15660 17684 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 7837 15555 7895 15561
rect 7837 15521 7849 15555
rect 7883 15552 7895 15555
rect 8110 15552 8116 15564
rect 7883 15524 8116 15552
rect 7883 15521 7895 15524
rect 7837 15515 7895 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 11514 15552 11520 15564
rect 11475 15524 11520 15552
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 14550 15552 14556 15564
rect 14511 15524 14556 15552
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15484 2927 15487
rect 4338 15484 4344 15496
rect 2915 15456 4344 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 4338 15444 4344 15456
rect 4396 15444 4402 15496
rect 5166 15484 5172 15496
rect 5127 15456 5172 15484
rect 5166 15444 5172 15456
rect 5224 15444 5230 15496
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7392 15456 7757 15484
rect 7282 15416 7288 15428
rect 6670 15388 7288 15416
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 7392 15360 7420 15456
rect 7745 15453 7757 15456
rect 7791 15453 7803 15487
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 7745 15447 7803 15453
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 10008 15456 10241 15484
rect 10008 15444 10014 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 10778 15484 10784 15496
rect 10459 15456 10784 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 14458 15484 14464 15496
rect 14419 15456 14464 15484
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 15378 15484 15384 15496
rect 15339 15456 15384 15484
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 15838 15484 15844 15496
rect 15611 15456 15844 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16022 15484 16028 15496
rect 15983 15456 16028 15484
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15484 16911 15487
rect 16942 15484 16948 15496
rect 16899 15456 16948 15484
rect 16899 15453 16911 15456
rect 16853 15447 16911 15453
rect 16942 15444 16948 15456
rect 17000 15484 17006 15496
rect 17494 15484 17500 15496
rect 17000 15456 17500 15484
rect 17000 15444 17006 15456
rect 17494 15444 17500 15456
rect 17552 15444 17558 15496
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 18288 15456 18337 15484
rect 18288 15444 18294 15456
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 18472 15456 18517 15484
rect 18472 15444 18478 15456
rect 11793 15419 11851 15425
rect 11793 15385 11805 15419
rect 11839 15385 11851 15419
rect 13354 15416 13360 15428
rect 13018 15388 13360 15416
rect 11793 15379 11851 15385
rect 3237 15351 3295 15357
rect 3237 15317 3249 15351
rect 3283 15348 3295 15351
rect 5258 15348 5264 15360
rect 3283 15320 5264 15348
rect 3283 15317 3295 15320
rect 3237 15311 3295 15317
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 7374 15348 7380 15360
rect 6963 15320 7380 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 11808 15348 11836 15379
rect 13354 15376 13360 15388
rect 13412 15376 13418 15428
rect 17126 15376 17132 15428
rect 17184 15416 17190 15428
rect 18141 15419 18199 15425
rect 18141 15416 18153 15419
rect 17184 15388 18153 15416
rect 17184 15376 17190 15388
rect 18141 15385 18153 15388
rect 18187 15385 18199 15419
rect 18141 15379 18199 15385
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 11808 15320 14105 15348
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 15194 15348 15200 15360
rect 15155 15320 15200 15348
rect 14093 15311 14151 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 16209 15351 16267 15357
rect 16209 15317 16221 15351
rect 16255 15348 16267 15351
rect 16574 15348 16580 15360
rect 16255 15320 16580 15348
rect 16255 15317 16267 15320
rect 16209 15311 16267 15317
rect 16574 15308 16580 15320
rect 16632 15348 16638 15360
rect 16758 15348 16764 15360
rect 16632 15320 16764 15348
rect 16632 15308 16638 15320
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 17589 15351 17647 15357
rect 17589 15317 17601 15351
rect 17635 15348 17647 15351
rect 17954 15348 17960 15360
rect 17635 15320 17960 15348
rect 17635 15317 17647 15320
rect 17589 15311 17647 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 1104 15258 19412 15280
rect 1104 15206 7052 15258
rect 7104 15206 7116 15258
rect 7168 15206 7180 15258
rect 7232 15206 7244 15258
rect 7296 15206 7308 15258
rect 7360 15206 13155 15258
rect 13207 15206 13219 15258
rect 13271 15206 13283 15258
rect 13335 15206 13347 15258
rect 13399 15206 13411 15258
rect 13463 15206 19412 15258
rect 1104 15184 19412 15206
rect 6914 15144 6920 15156
rect 6875 15116 6920 15144
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 12805 15147 12863 15153
rect 12805 15113 12817 15147
rect 12851 15144 12863 15147
rect 14458 15144 14464 15156
rect 12851 15116 14464 15144
rect 12851 15113 12863 15116
rect 12805 15107 12863 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 16574 15104 16580 15156
rect 16632 15144 16638 15156
rect 16942 15144 16948 15156
rect 16632 15116 16948 15144
rect 16632 15104 16638 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17310 15104 17316 15156
rect 17368 15104 17374 15156
rect 18414 15144 18420 15156
rect 18375 15116 18420 15144
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 6362 15036 6368 15088
rect 6420 15076 6426 15088
rect 6420 15048 7788 15076
rect 6420 15036 6426 15048
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 3878 15008 3884 15020
rect 2004 14980 3884 15008
rect 2004 14968 2010 14980
rect 3878 14968 3884 14980
rect 3936 15008 3942 15020
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 3936 14980 4629 15008
rect 3936 14968 3942 14980
rect 4617 14977 4629 14980
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 5261 15011 5319 15017
rect 5261 14977 5273 15011
rect 5307 15008 5319 15011
rect 6822 15008 6828 15020
rect 5307 14980 6828 15008
rect 5307 14977 5319 14980
rect 5261 14971 5319 14977
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 7101 15011 7159 15017
rect 7101 14977 7113 15011
rect 7147 14977 7159 15011
rect 7101 14971 7159 14977
rect 7285 15011 7343 15017
rect 7285 14977 7297 15011
rect 7331 15008 7343 15011
rect 7374 15008 7380 15020
rect 7331 14980 7380 15008
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 4522 14804 4528 14816
rect 4483 14776 4528 14804
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 7116 14804 7144 14971
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 7760 15017 7788 15048
rect 9030 15036 9036 15088
rect 9088 15036 9094 15088
rect 11514 15036 11520 15088
rect 11572 15076 11578 15088
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 11572 15048 11897 15076
rect 11572 15036 11578 15048
rect 11885 15045 11897 15048
rect 11931 15045 11943 15079
rect 11885 15039 11943 15045
rect 12069 15079 12127 15085
rect 12069 15045 12081 15079
rect 12115 15076 12127 15079
rect 13078 15076 13084 15088
rect 12115 15048 13084 15076
rect 12115 15045 12127 15048
rect 12069 15039 12127 15045
rect 13078 15036 13084 15048
rect 13136 15076 13142 15088
rect 13357 15079 13415 15085
rect 13357 15076 13369 15079
rect 13136 15048 13369 15076
rect 13136 15036 13142 15048
rect 13357 15045 13369 15048
rect 13403 15045 13415 15079
rect 15102 15076 15108 15088
rect 13357 15039 13415 15045
rect 14016 15048 15108 15076
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 10137 15011 10195 15017
rect 10137 15008 10149 15011
rect 10008 14980 10149 15008
rect 10008 14968 10014 14980
rect 10137 14977 10149 14980
rect 10183 14977 10195 15011
rect 10137 14971 10195 14977
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 11146 15008 11152 15020
rect 10367 14980 11152 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 14977 12679 15011
rect 12621 14971 12679 14977
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 15008 12863 15011
rect 14016 15008 14044 15048
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 15654 15076 15660 15088
rect 15304 15048 15660 15076
rect 12851 15006 13308 15008
rect 13464 15006 14044 15008
rect 12851 14980 14044 15006
rect 12851 14977 12863 14980
rect 13280 14978 13492 14980
rect 12805 14971 12863 14977
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 9214 14940 9220 14952
rect 8067 14912 9220 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 9214 14900 9220 14912
rect 9272 14900 9278 14952
rect 12636 14940 12664 14971
rect 14090 14968 14096 15020
rect 14148 15008 14154 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 14148 14980 14289 15008
rect 14148 14968 14154 14980
rect 14277 14977 14289 14980
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14461 15011 14519 15017
rect 14461 14977 14473 15011
rect 14507 15008 14519 15011
rect 15194 15008 15200 15020
rect 14507 14980 15200 15008
rect 14507 14977 14519 14980
rect 14461 14971 14519 14977
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 14108 14940 14136 14968
rect 12636 14912 14136 14940
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 15304 14940 15332 15048
rect 15654 15036 15660 15048
rect 15712 15076 15718 15088
rect 17328 15076 17356 15104
rect 15712 15048 17356 15076
rect 15712 15036 15718 15048
rect 17954 15036 17960 15088
rect 18012 15036 18018 15088
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 15838 15008 15844 15020
rect 15427 14980 15844 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 15470 14940 15476 14952
rect 14415 14912 15332 14940
rect 15431 14912 15476 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 14200 14872 14228 14903
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 16942 14940 16948 14952
rect 16903 14912 16948 14940
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 14550 14872 14556 14884
rect 14200 14844 14556 14872
rect 14550 14832 14556 14844
rect 14608 14872 14614 14884
rect 15013 14875 15071 14881
rect 15013 14872 15025 14875
rect 14608 14844 15025 14872
rect 14608 14832 14614 14844
rect 15013 14841 15025 14844
rect 15059 14841 15071 14875
rect 15013 14835 15071 14841
rect 8110 14804 8116 14816
rect 7116 14776 8116 14804
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 9493 14807 9551 14813
rect 9493 14773 9505 14807
rect 9539 14804 9551 14807
rect 9674 14804 9680 14816
rect 9539 14776 9680 14804
rect 9539 14773 9551 14776
rect 9493 14767 9551 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 10229 14807 10287 14813
rect 10229 14773 10241 14807
rect 10275 14804 10287 14807
rect 10502 14804 10508 14816
rect 10275 14776 10508 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 13446 14804 13452 14816
rect 13407 14776 13452 14804
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13998 14804 14004 14816
rect 13959 14776 14004 14804
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 1104 14714 19412 14736
rect 1104 14662 4001 14714
rect 4053 14662 4065 14714
rect 4117 14662 4129 14714
rect 4181 14662 4193 14714
rect 4245 14662 4257 14714
rect 4309 14662 10104 14714
rect 10156 14662 10168 14714
rect 10220 14662 10232 14714
rect 10284 14662 10296 14714
rect 10348 14662 10360 14714
rect 10412 14662 16206 14714
rect 16258 14662 16270 14714
rect 16322 14662 16334 14714
rect 16386 14662 16398 14714
rect 16450 14662 16462 14714
rect 16514 14662 19412 14714
rect 1104 14640 19412 14662
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 6089 14603 6147 14609
rect 6089 14600 6101 14603
rect 5132 14572 6101 14600
rect 5132 14560 5138 14572
rect 6089 14569 6101 14572
rect 6135 14569 6147 14603
rect 6089 14563 6147 14569
rect 2685 14467 2743 14473
rect 2685 14433 2697 14467
rect 2731 14464 2743 14467
rect 2731 14436 3740 14464
rect 2731 14433 2743 14436
rect 2685 14427 2743 14433
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 1946 14396 1952 14408
rect 1903 14368 1952 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14396 2835 14399
rect 3602 14396 3608 14408
rect 2823 14368 3608 14396
rect 2823 14365 2835 14368
rect 2777 14359 2835 14365
rect 1765 14331 1823 14337
rect 1765 14297 1777 14331
rect 1811 14328 1823 14331
rect 2130 14328 2136 14340
rect 1811 14300 2136 14328
rect 1811 14297 1823 14300
rect 1765 14291 1823 14297
rect 2130 14288 2136 14300
rect 2188 14288 2194 14340
rect 2608 14328 2636 14359
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 3712 14396 3740 14436
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 5166 14464 5172 14476
rect 3844 14436 5172 14464
rect 3844 14424 3850 14436
rect 5166 14424 5172 14436
rect 5224 14464 5230 14476
rect 5537 14467 5595 14473
rect 5537 14464 5549 14467
rect 5224 14436 5549 14464
rect 5224 14424 5230 14436
rect 5537 14433 5549 14436
rect 5583 14433 5595 14467
rect 6104 14464 6132 14563
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 6917 14603 6975 14609
rect 6917 14600 6929 14603
rect 6420 14572 6929 14600
rect 6420 14560 6426 14572
rect 6917 14569 6929 14572
rect 6963 14569 6975 14603
rect 6917 14563 6975 14569
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 7524 14572 7573 14600
rect 7524 14560 7530 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 9030 14600 9036 14612
rect 8991 14572 9036 14600
rect 7561 14563 7619 14569
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 14350 14603 14408 14609
rect 14350 14600 14362 14603
rect 14056 14572 14362 14600
rect 14056 14560 14062 14572
rect 14350 14569 14362 14572
rect 14396 14569 14408 14603
rect 15838 14600 15844 14612
rect 15799 14572 15844 14600
rect 14350 14563 14408 14569
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 16669 14603 16727 14609
rect 16669 14569 16681 14603
rect 16715 14600 16727 14603
rect 16942 14600 16948 14612
rect 16715 14572 16948 14600
rect 16715 14569 16727 14572
rect 16669 14563 16727 14569
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 16850 14492 16856 14544
rect 16908 14532 16914 14544
rect 17957 14535 18015 14541
rect 17957 14532 17969 14535
rect 16908 14504 17969 14532
rect 16908 14492 16914 14504
rect 17957 14501 17969 14504
rect 18003 14501 18015 14535
rect 17957 14495 18015 14501
rect 10318 14464 10324 14476
rect 6104 14436 7512 14464
rect 10279 14436 10324 14464
rect 5537 14427 5595 14433
rect 3712 14368 3924 14396
rect 3510 14328 3516 14340
rect 2608 14300 3516 14328
rect 3510 14288 3516 14300
rect 3568 14288 3574 14340
rect 1946 14220 1952 14272
rect 2004 14260 2010 14272
rect 2317 14263 2375 14269
rect 2317 14260 2329 14263
rect 2004 14232 2329 14260
rect 2004 14220 2010 14232
rect 2317 14229 2329 14232
rect 2363 14229 2375 14263
rect 2317 14223 2375 14229
rect 3694 14220 3700 14272
rect 3752 14260 3758 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3752 14232 3801 14260
rect 3752 14220 3758 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 3896 14260 3924 14368
rect 6178 14356 6184 14408
rect 6236 14396 6242 14408
rect 6273 14399 6331 14405
rect 6273 14396 6285 14399
rect 6236 14368 6285 14396
rect 6236 14356 6242 14368
rect 6273 14365 6285 14368
rect 6319 14365 6331 14399
rect 6822 14396 6828 14408
rect 6783 14368 6828 14396
rect 6273 14359 6331 14365
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 7484 14405 7512 14436
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13504 14436 14105 14464
rect 13504 14424 13510 14436
rect 14093 14433 14105 14436
rect 14139 14464 14151 14467
rect 16666 14464 16672 14476
rect 14139 14436 16672 14464
rect 14139 14433 14151 14436
rect 14093 14427 14151 14433
rect 16666 14424 16672 14436
rect 16724 14424 16730 14476
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 16816 14436 16957 14464
rect 16816 14424 16822 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 17126 14464 17132 14476
rect 17087 14436 17132 14464
rect 16945 14427 17003 14433
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 18230 14464 18236 14476
rect 18143 14436 18236 14464
rect 18230 14424 18236 14436
rect 18288 14464 18294 14476
rect 18690 14464 18696 14476
rect 18288 14436 18696 14464
rect 18288 14424 18294 14436
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14365 7527 14399
rect 9122 14396 9128 14408
rect 9083 14368 9128 14396
rect 7469 14359 7527 14365
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 10502 14396 10508 14408
rect 10459 14368 10508 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 11425 14399 11483 14405
rect 11425 14365 11437 14399
rect 11471 14365 11483 14399
rect 11425 14359 11483 14365
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14396 12403 14399
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 12391 14368 13553 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 13541 14365 13553 14368
rect 13587 14396 13599 14399
rect 13998 14396 14004 14408
rect 13587 14368 14004 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 4522 14288 4528 14340
rect 4580 14288 4586 14340
rect 5258 14328 5264 14340
rect 5219 14300 5264 14328
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 9140 14328 9168 14356
rect 11440 14328 11468 14359
rect 13998 14356 14004 14368
rect 14056 14356 14062 14408
rect 16850 14396 16856 14408
rect 16811 14368 16856 14396
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14396 17095 14399
rect 17310 14396 17316 14408
rect 17083 14368 17316 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18414 14396 18420 14408
rect 18371 14368 18420 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 9140 14300 12204 14328
rect 4338 14260 4344 14272
rect 3896 14232 4344 14260
rect 3789 14223 3847 14229
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 10781 14263 10839 14269
rect 10781 14229 10793 14263
rect 10827 14260 10839 14263
rect 11422 14260 11428 14272
rect 10827 14232 11428 14260
rect 10827 14229 10839 14232
rect 10781 14223 10839 14229
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 11517 14263 11575 14269
rect 11517 14229 11529 14263
rect 11563 14260 11575 14263
rect 11882 14260 11888 14272
rect 11563 14232 11888 14260
rect 11563 14229 11575 14232
rect 11517 14223 11575 14229
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 12176 14269 12204 14300
rect 15378 14288 15384 14340
rect 15436 14288 15442 14340
rect 12161 14263 12219 14269
rect 12161 14229 12173 14263
rect 12207 14229 12219 14263
rect 12161 14223 12219 14229
rect 13357 14263 13415 14269
rect 13357 14229 13369 14263
rect 13403 14260 13415 14263
rect 13630 14260 13636 14272
rect 13403 14232 13636 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 1104 14170 19412 14192
rect 1104 14118 7052 14170
rect 7104 14118 7116 14170
rect 7168 14118 7180 14170
rect 7232 14118 7244 14170
rect 7296 14118 7308 14170
rect 7360 14118 13155 14170
rect 13207 14118 13219 14170
rect 13271 14118 13283 14170
rect 13335 14118 13347 14170
rect 13399 14118 13411 14170
rect 13463 14118 19412 14170
rect 1104 14096 19412 14118
rect 3786 14056 3792 14068
rect 1412 14028 3792 14056
rect 1412 13929 1440 14028
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 3878 14016 3884 14068
rect 3936 14056 3942 14068
rect 4617 14059 4675 14065
rect 4617 14056 4629 14059
rect 3936 14028 4629 14056
rect 3936 14016 3942 14028
rect 4617 14025 4629 14028
rect 4663 14025 4675 14059
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 4617 14019 4675 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 15013 14059 15071 14065
rect 15013 14025 15025 14059
rect 15059 14056 15071 14059
rect 15102 14056 15108 14068
rect 15059 14028 15108 14056
rect 15059 14025 15071 14028
rect 15013 14019 15071 14025
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 16574 14056 16580 14068
rect 15887 14028 16580 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 16853 14059 16911 14065
rect 16853 14025 16865 14059
rect 16899 14056 16911 14059
rect 17954 14056 17960 14068
rect 16899 14028 17960 14056
rect 16899 14025 16911 14028
rect 16853 14019 16911 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 1946 13988 1952 14000
rect 1719 13960 1952 13988
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 1946 13948 1952 13960
rect 2004 13948 2010 14000
rect 2130 13948 2136 14000
rect 2188 13948 2194 14000
rect 3602 13988 3608 14000
rect 3563 13960 3608 13988
rect 3602 13948 3608 13960
rect 3660 13948 3666 14000
rect 8938 13988 8944 14000
rect 7866 13960 8944 13988
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 11146 13988 11152 14000
rect 10520 13960 11152 13988
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 3694 13880 3700 13932
rect 3752 13920 3758 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3752 13892 3801 13920
rect 3752 13880 3758 13892
rect 3789 13889 3801 13892
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13920 4859 13923
rect 6178 13920 6184 13932
rect 4847 13892 6184 13920
rect 4847 13889 4859 13892
rect 4801 13883 4859 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 6362 13920 6368 13932
rect 6323 13892 6368 13920
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 9364 13892 9413 13920
rect 9364 13880 9370 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 10318 13920 10324 13932
rect 9401 13883 9459 13889
rect 9784 13892 10324 13920
rect 3142 13852 3148 13864
rect 3055 13824 3148 13852
rect 3142 13812 3148 13824
rect 3200 13852 3206 13864
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 3200 13824 3985 13852
rect 3200 13812 3206 13824
rect 3973 13821 3985 13824
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13852 9551 13855
rect 9674 13852 9680 13864
rect 9539 13824 9680 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 9784 13861 9812 13892
rect 10318 13880 10324 13892
rect 10376 13920 10382 13932
rect 10520 13929 10548 13960
rect 11146 13948 11152 13960
rect 11204 13948 11210 14000
rect 11422 13948 11428 14000
rect 11480 13988 11486 14000
rect 11793 13991 11851 13997
rect 11793 13988 11805 13991
rect 11480 13960 11805 13988
rect 11480 13948 11486 13960
rect 11793 13957 11805 13960
rect 11839 13957 11851 13991
rect 11793 13951 11851 13957
rect 11882 13948 11888 14000
rect 11940 13988 11946 14000
rect 11940 13960 12282 13988
rect 11940 13948 11946 13960
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 13725 13991 13783 13997
rect 13725 13988 13737 13991
rect 13136 13960 13737 13988
rect 13136 13948 13142 13960
rect 13725 13957 13737 13960
rect 13771 13957 13783 13991
rect 13725 13951 13783 13957
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 10376 13892 10425 13920
rect 10376 13880 10382 13892
rect 10413 13889 10425 13892
rect 10459 13889 10471 13923
rect 10413 13883 10471 13889
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 10962 13920 10968 13932
rect 10643 13892 10968 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11514 13920 11520 13932
rect 11112 13892 11520 13920
rect 11112 13880 11118 13892
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14182 13920 14188 13932
rect 13955 13892 14188 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13889 15715 13923
rect 15657 13883 15715 13889
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 17034 13920 17040 13932
rect 16715 13892 17040 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 10229 13855 10287 13861
rect 10229 13852 10241 13855
rect 9916 13824 10241 13852
rect 9916 13812 9922 13824
rect 10229 13821 10241 13824
rect 10275 13821 10287 13855
rect 10229 13815 10287 13821
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 10744 13824 10789 13852
rect 10744 13812 10750 13824
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14826 13852 14832 13864
rect 14056 13824 14832 13852
rect 14056 13812 14062 13824
rect 14826 13812 14832 13824
rect 14884 13852 14890 13864
rect 15672 13852 15700 13883
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 14884 13824 15700 13852
rect 14884 13812 14890 13824
rect 6086 13676 6092 13728
rect 6144 13716 6150 13728
rect 6622 13719 6680 13725
rect 6622 13716 6634 13719
rect 6144 13688 6634 13716
rect 6144 13676 6150 13688
rect 6622 13685 6634 13688
rect 6668 13685 6680 13719
rect 6622 13679 6680 13685
rect 13265 13719 13323 13725
rect 13265 13685 13277 13719
rect 13311 13716 13323 13719
rect 13538 13716 13544 13728
rect 13311 13688 13544 13716
rect 13311 13685 13323 13688
rect 13265 13679 13323 13685
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 1104 13626 19412 13648
rect 1104 13574 4001 13626
rect 4053 13574 4065 13626
rect 4117 13574 4129 13626
rect 4181 13574 4193 13626
rect 4245 13574 4257 13626
rect 4309 13574 10104 13626
rect 10156 13574 10168 13626
rect 10220 13574 10232 13626
rect 10284 13574 10296 13626
rect 10348 13574 10360 13626
rect 10412 13574 16206 13626
rect 16258 13574 16270 13626
rect 16322 13574 16334 13626
rect 16386 13574 16398 13626
rect 16450 13574 16462 13626
rect 16514 13574 19412 13626
rect 1104 13552 19412 13574
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 2498 13512 2504 13524
rect 2271 13484 2504 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6733 13515 6791 13521
rect 6733 13481 6745 13515
rect 6779 13512 6791 13515
rect 6822 13512 6828 13524
rect 6779 13484 6828 13512
rect 6779 13481 6791 13484
rect 6733 13475 6791 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10686 13512 10692 13524
rect 10091 13484 10692 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 14185 13515 14243 13521
rect 11020 13484 12434 13512
rect 11020 13472 11026 13484
rect 7653 13447 7711 13453
rect 7653 13444 7665 13447
rect 5276 13416 7665 13444
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13376 2743 13379
rect 3694 13376 3700 13388
rect 2731 13348 3700 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 3694 13336 3700 13348
rect 3752 13336 3758 13388
rect 4430 13376 4436 13388
rect 3804 13348 4436 13376
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13308 2651 13311
rect 3142 13308 3148 13320
rect 2639 13280 3148 13308
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3510 13268 3516 13320
rect 3568 13308 3574 13320
rect 3804 13317 3832 13348
rect 4430 13336 4436 13348
rect 4488 13336 4494 13388
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3568 13280 3801 13308
rect 3568 13268 3574 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4614 13308 4620 13320
rect 4019 13280 4620 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4614 13268 4620 13280
rect 4672 13308 4678 13320
rect 5276 13308 5304 13416
rect 7653 13413 7665 13416
rect 7699 13413 7711 13447
rect 7653 13407 7711 13413
rect 11330 13404 11336 13456
rect 11388 13404 11394 13456
rect 5902 13376 5908 13388
rect 5863 13348 5908 13376
rect 5902 13336 5908 13348
rect 5960 13336 5966 13388
rect 11348 13376 11376 13404
rect 11532 13385 11560 13484
rect 12406 13444 12434 13484
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 15378 13512 15384 13524
rect 14231 13484 15384 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 18690 13512 18696 13524
rect 18651 13484 18696 13512
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 12529 13447 12587 13453
rect 12529 13444 12541 13447
rect 12406 13416 12541 13444
rect 12529 13413 12541 13416
rect 12575 13413 12587 13447
rect 12529 13407 12587 13413
rect 11425 13379 11483 13385
rect 11425 13376 11437 13379
rect 11348 13348 11437 13376
rect 11425 13345 11437 13348
rect 11471 13345 11483 13379
rect 11425 13339 11483 13345
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 13446 13336 13452 13388
rect 13504 13376 13510 13388
rect 14734 13376 14740 13388
rect 13504 13348 14740 13376
rect 13504 13336 13510 13348
rect 14734 13336 14740 13348
rect 14792 13376 14798 13388
rect 16022 13376 16028 13388
rect 14792 13348 14872 13376
rect 15983 13348 16028 13376
rect 14792 13336 14798 13348
rect 4672 13280 5304 13308
rect 5813 13311 5871 13317
rect 4672 13268 4678 13280
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 7466 13308 7472 13320
rect 5859 13280 7472 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 9306 13308 9312 13320
rect 8444 13280 9312 13308
rect 8444 13268 8450 13280
rect 9306 13268 9312 13280
rect 9364 13308 9370 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9364 13280 9689 13308
rect 9364 13268 9370 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 9861 13311 9919 13317
rect 9861 13308 9873 13311
rect 9824 13280 9873 13308
rect 9824 13268 9830 13280
rect 9861 13277 9873 13280
rect 9907 13277 9919 13311
rect 9861 13271 9919 13277
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 10560 13280 11345 13308
rect 10560 13268 10566 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 11664 13280 11709 13308
rect 11664 13268 11670 13280
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 14844 13317 14872 13348
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16666 13336 16672 13388
rect 16724 13376 16730 13388
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 16724 13348 16957 13376
rect 16724 13336 16730 13348
rect 16945 13345 16957 13348
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13688 13280 14105 13308
rect 13688 13268 13694 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13277 14887 13311
rect 16114 13308 16120 13320
rect 16075 13280 16120 13308
rect 14829 13271 14887 13277
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 6825 13243 6883 13249
rect 6825 13209 6837 13243
rect 6871 13240 6883 13243
rect 6914 13240 6920 13252
rect 6871 13212 6920 13240
rect 6871 13209 6883 13212
rect 6825 13203 6883 13209
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 7834 13240 7840 13252
rect 7795 13212 7840 13240
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 12713 13243 12771 13249
rect 12713 13209 12725 13243
rect 12759 13240 12771 13243
rect 13998 13240 14004 13252
rect 12759 13212 14004 13240
rect 12759 13209 12771 13212
rect 12713 13203 12771 13209
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 17221 13243 17279 13249
rect 17221 13240 17233 13243
rect 16500 13212 17233 13240
rect 2590 13132 2596 13184
rect 2648 13172 2654 13184
rect 3881 13175 3939 13181
rect 3881 13172 3893 13175
rect 2648 13144 3893 13172
rect 2648 13132 2654 13144
rect 3881 13141 3893 13144
rect 3927 13141 3939 13175
rect 11146 13172 11152 13184
rect 11107 13144 11152 13172
rect 3881 13135 3939 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 13964 13144 14933 13172
rect 13964 13132 13970 13144
rect 14921 13141 14933 13144
rect 14967 13172 14979 13175
rect 15102 13172 15108 13184
rect 14967 13144 15108 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 16500 13181 16528 13212
rect 17221 13209 17233 13212
rect 17267 13209 17279 13243
rect 18506 13240 18512 13252
rect 18446 13212 18512 13240
rect 17221 13203 17279 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 16485 13175 16543 13181
rect 16485 13141 16497 13175
rect 16531 13141 16543 13175
rect 16485 13135 16543 13141
rect 1104 13082 19412 13104
rect 1104 13030 7052 13082
rect 7104 13030 7116 13082
rect 7168 13030 7180 13082
rect 7232 13030 7244 13082
rect 7296 13030 7308 13082
rect 7360 13030 13155 13082
rect 13207 13030 13219 13082
rect 13271 13030 13283 13082
rect 13335 13030 13347 13082
rect 13399 13030 13411 13082
rect 13463 13030 19412 13082
rect 1104 13008 19412 13030
rect 4893 12971 4951 12977
rect 4893 12937 4905 12971
rect 4939 12968 4951 12971
rect 5534 12968 5540 12980
rect 4939 12940 5540 12968
rect 4939 12937 4951 12940
rect 4893 12931 4951 12937
rect 5534 12928 5540 12940
rect 5592 12968 5598 12980
rect 6730 12968 6736 12980
rect 5592 12940 6736 12968
rect 5592 12928 5598 12940
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 7466 12968 7472 12980
rect 7427 12940 7472 12968
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 8938 12968 8944 12980
rect 8899 12940 8944 12968
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 11664 12940 13369 12968
rect 11664 12928 11670 12940
rect 13357 12937 13369 12940
rect 13403 12937 13415 12971
rect 15654 12968 15660 12980
rect 15615 12940 15660 12968
rect 13357 12931 13415 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 16172 12940 17785 12968
rect 16172 12928 16178 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 18506 12968 18512 12980
rect 18467 12940 18512 12968
rect 17773 12931 17831 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 7650 12900 7656 12912
rect 7392 12872 7656 12900
rect 2590 12832 2596 12844
rect 2551 12804 2596 12832
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3936 12804 3985 12832
rect 3936 12792 3942 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 4982 12832 4988 12844
rect 4943 12804 4988 12832
rect 3973 12795 4031 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 6546 12832 6552 12844
rect 5960 12804 6552 12832
rect 5960 12792 5966 12804
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 7392 12841 7420 12872
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 7834 12860 7840 12912
rect 7892 12900 7898 12912
rect 8297 12903 8355 12909
rect 8297 12900 8309 12903
rect 7892 12872 8309 12900
rect 7892 12860 7898 12872
rect 8297 12869 8309 12872
rect 8343 12900 8355 12903
rect 9953 12903 10011 12909
rect 9953 12900 9965 12903
rect 8343 12872 9965 12900
rect 8343 12869 8355 12872
rect 8297 12863 8355 12869
rect 9953 12869 9965 12872
rect 9999 12900 10011 12903
rect 13906 12900 13912 12912
rect 9999 12872 13912 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 13998 12860 14004 12912
rect 14056 12900 14062 12912
rect 15565 12903 15623 12909
rect 15565 12900 15577 12903
rect 14056 12872 15577 12900
rect 14056 12860 14062 12872
rect 15565 12869 15577 12872
rect 15611 12869 15623 12903
rect 15565 12863 15623 12869
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6687 12804 7389 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 7607 12804 8125 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 8113 12801 8125 12804
rect 8159 12832 8171 12835
rect 8202 12832 8208 12844
rect 8159 12804 8208 12832
rect 8159 12801 8171 12804
rect 8113 12795 8171 12801
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 8846 12832 8852 12844
rect 8807 12804 8852 12832
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 12710 12832 12716 12844
rect 12671 12804 12716 12832
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 13538 12832 13544 12844
rect 12820 12804 13544 12832
rect 2498 12764 2504 12776
rect 2459 12736 2504 12764
rect 2498 12724 2504 12736
rect 2556 12724 2562 12776
rect 6730 12764 6736 12776
rect 6691 12736 6736 12764
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 9769 12767 9827 12773
rect 6871 12736 7420 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7392 12708 7420 12736
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 9950 12764 9956 12776
rect 9815 12736 9956 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 9950 12724 9956 12736
rect 10008 12724 10014 12776
rect 10502 12724 10508 12776
rect 10560 12764 10566 12776
rect 12820 12773 12848 12804
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 14734 12832 14740 12844
rect 14695 12804 14740 12832
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 15160 12804 17141 12832
rect 15160 12792 15166 12804
rect 17129 12801 17141 12804
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17773 12835 17831 12841
rect 17773 12832 17785 12835
rect 17368 12804 17785 12832
rect 17368 12792 17374 12804
rect 17773 12801 17785 12804
rect 17819 12801 17831 12835
rect 17954 12832 17960 12844
rect 17915 12804 17960 12832
rect 17773 12795 17831 12801
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 10560 12736 12357 12764
rect 10560 12724 10566 12736
rect 12345 12733 12357 12736
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 13722 12764 13728 12776
rect 13683 12736 13728 12764
rect 12805 12727 12863 12733
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 18432 12764 18460 12795
rect 16816 12736 18460 12764
rect 16816 12724 16822 12736
rect 2958 12696 2964 12708
rect 2919 12668 2964 12696
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 4982 12656 4988 12708
rect 5040 12696 5046 12708
rect 5040 12668 6500 12696
rect 5040 12656 5046 12668
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4522 12628 4528 12640
rect 4111 12600 4528 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 6362 12628 6368 12640
rect 6323 12600 6368 12628
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 6472 12628 6500 12668
rect 7374 12656 7380 12708
rect 7432 12656 7438 12708
rect 12406 12668 14412 12696
rect 12406 12628 12434 12668
rect 14384 12640 14412 12668
rect 6472 12600 12434 12628
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 14921 12631 14979 12637
rect 14921 12628 14933 12631
rect 14424 12600 14933 12628
rect 14424 12588 14430 12600
rect 14921 12597 14933 12600
rect 14967 12597 14979 12631
rect 14921 12591 14979 12597
rect 1104 12538 19412 12560
rect 1104 12486 4001 12538
rect 4053 12486 4065 12538
rect 4117 12486 4129 12538
rect 4181 12486 4193 12538
rect 4245 12486 4257 12538
rect 4309 12486 10104 12538
rect 10156 12486 10168 12538
rect 10220 12486 10232 12538
rect 10284 12486 10296 12538
rect 10348 12486 10360 12538
rect 10412 12486 16206 12538
rect 16258 12486 16270 12538
rect 16322 12486 16334 12538
rect 16386 12486 16398 12538
rect 16450 12486 16462 12538
rect 16514 12486 19412 12538
rect 1104 12464 19412 12486
rect 6546 12384 6552 12436
rect 6604 12424 6610 12436
rect 6825 12427 6883 12433
rect 6825 12424 6837 12427
rect 6604 12396 6837 12424
rect 6604 12384 6610 12396
rect 6825 12393 6837 12396
rect 6871 12393 6883 12427
rect 11330 12424 11336 12436
rect 6825 12387 6883 12393
rect 10428 12396 11336 12424
rect 3786 12288 3792 12300
rect 3747 12260 3792 12288
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12288 7343 12291
rect 7374 12288 7380 12300
rect 7331 12260 7380 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7558 12220 7564 12232
rect 7239 12192 7564 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10428 12229 10456 12396
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 12621 12427 12679 12433
rect 12621 12393 12633 12427
rect 12667 12424 12679 12427
rect 12710 12424 12716 12436
rect 12667 12396 12716 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 12710 12384 12716 12396
rect 12768 12424 12774 12436
rect 13722 12424 13728 12436
rect 12768 12396 13728 12424
rect 12768 12384 12774 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 11146 12288 11152 12300
rect 11107 12260 11152 12288
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12288 14611 12291
rect 14734 12288 14740 12300
rect 14599 12260 14740 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 16393 12291 16451 12297
rect 16393 12288 16405 12291
rect 15712 12260 16405 12288
rect 15712 12248 15718 12260
rect 16393 12257 16405 12260
rect 16439 12257 16451 12291
rect 16393 12251 16451 12257
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10008 12192 10241 12220
rect 10008 12180 10014 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 2958 12112 2964 12164
rect 3016 12152 3022 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 3016 12124 4077 12152
rect 3016 12112 3022 12124
rect 4065 12121 4077 12124
rect 4111 12121 4123 12155
rect 4065 12115 4123 12121
rect 4522 12112 4528 12164
rect 4580 12112 4586 12164
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7834 12152 7840 12164
rect 6972 12124 7840 12152
rect 6972 12112 6978 12124
rect 7834 12112 7840 12124
rect 7892 12112 7898 12164
rect 8018 12152 8024 12164
rect 7979 12124 8024 12152
rect 8018 12112 8024 12124
rect 8076 12112 8082 12164
rect 10888 12152 10916 12183
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14056 12192 14841 12220
rect 14056 12180 14062 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 16206 12220 16212 12232
rect 16167 12192 16212 12220
rect 14829 12183 14887 12189
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12220 16543 12223
rect 17862 12220 17868 12232
rect 16531 12192 17868 12220
rect 16531 12189 16543 12192
rect 16485 12183 16543 12189
rect 11054 12152 11060 12164
rect 10888 12124 11060 12152
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 11882 12112 11888 12164
rect 11940 12112 11946 12164
rect 16316 12152 16344 12183
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 17954 12152 17960 12164
rect 16316 12124 17960 12152
rect 17954 12112 17960 12124
rect 18012 12112 18018 12164
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 4764 12056 5549 12084
rect 4764 12044 4770 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 10321 12087 10379 12093
rect 10321 12053 10333 12087
rect 10367 12084 10379 12087
rect 10594 12084 10600 12096
rect 10367 12056 10600 12084
rect 10367 12053 10379 12056
rect 10321 12047 10379 12053
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15988 12056 16037 12084
rect 15988 12044 15994 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 1104 11994 19412 12016
rect 1104 11942 7052 11994
rect 7104 11942 7116 11994
rect 7168 11942 7180 11994
rect 7232 11942 7244 11994
rect 7296 11942 7308 11994
rect 7360 11942 13155 11994
rect 13207 11942 13219 11994
rect 13271 11942 13283 11994
rect 13335 11942 13347 11994
rect 13399 11942 13411 11994
rect 13463 11942 19412 11994
rect 1104 11920 19412 11942
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11880 6975 11883
rect 7466 11880 7472 11892
rect 6963 11852 7472 11880
rect 6963 11849 6975 11852
rect 6917 11843 6975 11849
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 8386 11880 8392 11892
rect 8347 11852 8392 11880
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 9692 11852 10701 11880
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 4525 11815 4583 11821
rect 4525 11812 4537 11815
rect 4396 11784 4537 11812
rect 4396 11772 4402 11784
rect 4525 11781 4537 11784
rect 4571 11781 4583 11815
rect 4525 11775 4583 11781
rect 4709 11815 4767 11821
rect 4709 11781 4721 11815
rect 4755 11812 4767 11815
rect 4982 11812 4988 11824
rect 4755 11784 4988 11812
rect 4755 11781 4767 11784
rect 4709 11775 4767 11781
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 9692 11812 9720 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11940 11852 11989 11880
rect 11940 11840 11946 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 11977 11843 12035 11849
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 14734 11880 14740 11892
rect 14507 11852 14740 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 9858 11812 9864 11824
rect 9430 11784 9720 11812
rect 9819 11784 9864 11812
rect 9858 11772 9864 11784
rect 9916 11772 9922 11824
rect 13541 11815 13599 11821
rect 13541 11781 13553 11815
rect 13587 11812 13599 11815
rect 18138 11812 18144 11824
rect 13587 11784 18144 11812
rect 13587 11781 13599 11784
rect 13541 11775 13599 11781
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 3418 11744 3424 11756
rect 2547 11716 3424 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 7374 11744 7380 11756
rect 7147 11716 7380 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 5828 11608 5856 11707
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 10827 11716 11897 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11885 11713 11897 11716
rect 11931 11744 11943 11747
rect 12342 11744 12348 11756
rect 11931 11716 12348 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 12710 11704 12716 11756
rect 12768 11744 12774 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 12768 11716 13369 11744
rect 12768 11704 12774 11716
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11744 13691 11747
rect 13998 11744 14004 11756
rect 13679 11716 14004 11744
rect 13679 11713 13691 11716
rect 13633 11707 13691 11713
rect 7282 11676 7288 11688
rect 7243 11648 7288 11676
rect 7282 11636 7288 11648
rect 7340 11676 7346 11688
rect 7558 11676 7564 11688
rect 7340 11648 7564 11676
rect 7340 11636 7346 11648
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 11054 11676 11060 11688
rect 10183 11648 11060 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 13372 11676 13400 11707
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14568 11753 14596 11784
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 14553 11747 14611 11753
rect 14553 11713 14565 11747
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 14292 11676 14320 11707
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 14884 11716 15025 11744
rect 14884 11704 14890 11716
rect 15013 11713 15025 11716
rect 15059 11713 15071 11747
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15013 11707 15071 11713
rect 15212 11716 16681 11744
rect 13372 11648 14320 11676
rect 6454 11608 6460 11620
rect 5828 11580 6460 11608
rect 6454 11568 6460 11580
rect 6512 11608 6518 11620
rect 8846 11608 8852 11620
rect 6512 11580 8852 11608
rect 6512 11568 6518 11580
rect 8846 11568 8852 11580
rect 8904 11568 8910 11620
rect 12805 11611 12863 11617
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 14182 11608 14188 11620
rect 12851 11580 14188 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 15212 11617 15240 11716
rect 16669 11713 16681 11716
rect 16715 11744 16727 11747
rect 16758 11744 16764 11756
rect 16715 11716 16764 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 18012 11716 18061 11744
rect 18012 11704 18018 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 16206 11636 16212 11688
rect 16264 11676 16270 11688
rect 17681 11679 17739 11685
rect 17681 11676 17693 11679
rect 16264 11648 17693 11676
rect 16264 11636 16270 11648
rect 17681 11645 17693 11648
rect 17727 11645 17739 11679
rect 18141 11679 18199 11685
rect 18141 11676 18153 11679
rect 17681 11639 17739 11645
rect 18064 11648 18153 11676
rect 18064 11620 18092 11648
rect 18141 11645 18153 11648
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 15197 11611 15255 11617
rect 15197 11577 15209 11611
rect 15243 11577 15255 11611
rect 15197 11571 15255 11577
rect 18046 11568 18052 11620
rect 18104 11568 18110 11620
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2406 11540 2412 11552
rect 2367 11512 2412 11540
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 5718 11540 5724 11552
rect 5679 11512 5724 11540
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 14090 11540 14096 11552
rect 14051 11512 14096 11540
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16724 11512 16773 11540
rect 16724 11500 16730 11512
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 16761 11503 16819 11509
rect 1104 11450 19412 11472
rect 1104 11398 4001 11450
rect 4053 11398 4065 11450
rect 4117 11398 4129 11450
rect 4181 11398 4193 11450
rect 4245 11398 4257 11450
rect 4309 11398 10104 11450
rect 10156 11398 10168 11450
rect 10220 11398 10232 11450
rect 10284 11398 10296 11450
rect 10348 11398 10360 11450
rect 10412 11398 16206 11450
rect 16258 11398 16270 11450
rect 16322 11398 16334 11450
rect 16386 11398 16398 11450
rect 16450 11398 16462 11450
rect 16514 11398 19412 11450
rect 1104 11376 19412 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 6549 11339 6607 11345
rect 6549 11305 6561 11339
rect 6595 11336 6607 11339
rect 7282 11336 7288 11348
rect 6595 11308 7288 11336
rect 6595 11305 6607 11308
rect 6549 11299 6607 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 17862 11336 17868 11348
rect 17823 11308 17868 11336
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 7561 11271 7619 11277
rect 7561 11237 7573 11271
rect 7607 11268 7619 11271
rect 8294 11268 8300 11280
rect 7607 11240 8300 11268
rect 7607 11237 7619 11240
rect 7561 11231 7619 11237
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 6362 11200 6368 11212
rect 5123 11172 6368 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6972 11172 7113 11200
rect 6972 11160 6978 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 8076 11172 10149 11200
rect 8076 11160 8082 11172
rect 10137 11169 10149 11172
rect 10183 11200 10195 11203
rect 12618 11200 12624 11212
rect 10183 11172 12624 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 14090 11200 14096 11212
rect 14051 11172 14096 11200
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 16574 11200 16580 11212
rect 15703 11172 16580 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 17954 11200 17960 11212
rect 17451 11172 17960 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 17954 11160 17960 11172
rect 18012 11200 18018 11212
rect 18233 11203 18291 11209
rect 18233 11200 18245 11203
rect 18012 11172 18245 11200
rect 18012 11160 18018 11172
rect 18233 11169 18245 11172
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3694 11132 3700 11144
rect 3191 11104 3700 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3694 11092 3700 11104
rect 3752 11132 3758 11144
rect 4801 11135 4859 11141
rect 4801 11132 4813 11135
rect 3752 11104 4813 11132
rect 3752 11092 3758 11104
rect 4801 11101 4813 11104
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8846 11132 8852 11144
rect 8251 11104 8852 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 2406 11024 2412 11076
rect 2464 11024 2470 11076
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 2832 11036 2881 11064
rect 2832 11024 2838 11036
rect 2869 11033 2881 11036
rect 2915 11033 2927 11067
rect 2869 11027 2927 11033
rect 5718 11024 5724 11076
rect 5776 11024 5782 11076
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 7208 10996 7236 11095
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9582 11132 9588 11144
rect 9539 11104 9588 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9324 11064 9352 11095
rect 9582 11092 9588 11104
rect 9640 11132 9646 11144
rect 11698 11132 11704 11144
rect 9640 11104 11704 11132
rect 9640 11092 9646 11104
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 13044 11104 13185 11132
rect 13044 11092 13050 11104
rect 13173 11101 13185 11104
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11132 13323 11135
rect 13538 11132 13544 11144
rect 13311 11104 13544 11132
rect 13311 11101 13323 11104
rect 13265 11095 13323 11101
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 13630 11092 13636 11144
rect 13688 11132 13694 11144
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 13688 11104 14289 11132
rect 13688 11092 13694 11104
rect 14277 11101 14289 11104
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 15562 11132 15568 11144
rect 14507 11104 15568 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 9950 11064 9956 11076
rect 9324 11036 9956 11064
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 11885 11067 11943 11073
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 15838 11064 15844 11076
rect 11931 11036 15844 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 15930 11024 15936 11076
rect 15988 11064 15994 11076
rect 15988 11036 16033 11064
rect 15988 11024 15994 11036
rect 16666 11024 16672 11076
rect 16724 11024 16730 11076
rect 6696 10968 7236 10996
rect 6696 10956 6702 10968
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8113 10999 8171 11005
rect 8113 10996 8125 10999
rect 8076 10968 8125 10996
rect 8076 10956 8082 10968
rect 8113 10965 8125 10968
rect 8159 10965 8171 10999
rect 9306 10996 9312 11008
rect 9267 10968 9312 10996
rect 8113 10959 8171 10965
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12492 10968 12537 10996
rect 12492 10956 12498 10968
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 17310 10996 17316 11008
rect 15252 10968 17316 10996
rect 15252 10956 15258 10968
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 1104 10906 19412 10928
rect 1104 10854 7052 10906
rect 7104 10854 7116 10906
rect 7168 10854 7180 10906
rect 7232 10854 7244 10906
rect 7296 10854 7308 10906
rect 7360 10854 13155 10906
rect 13207 10854 13219 10906
rect 13271 10854 13283 10906
rect 13335 10854 13347 10906
rect 13399 10854 13411 10906
rect 13463 10854 19412 10906
rect 1104 10832 19412 10854
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 6638 10792 6644 10804
rect 5859 10764 6644 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 6825 10795 6883 10801
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 7374 10792 7380 10804
rect 6871 10764 7380 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 12710 10792 12716 10804
rect 12671 10764 12716 10792
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 16117 10795 16175 10801
rect 16117 10761 16129 10795
rect 16163 10761 16175 10795
rect 16117 10755 16175 10761
rect 5994 10724 6000 10736
rect 5644 10696 6000 10724
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 2958 10656 2964 10668
rect 2915 10628 2964 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3326 10656 3332 10668
rect 3099 10628 3332 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 5644 10665 5672 10696
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 8018 10724 8024 10736
rect 7866 10696 8024 10724
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 8294 10724 8300 10736
rect 8255 10696 8300 10724
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 13538 10684 13544 10736
rect 13596 10684 13602 10736
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 14185 10727 14243 10733
rect 14185 10724 14197 10727
rect 14148 10696 14197 10724
rect 14148 10684 14154 10696
rect 14185 10693 14197 10696
rect 14231 10693 14243 10727
rect 14185 10687 14243 10693
rect 15013 10727 15071 10733
rect 15013 10693 15025 10727
rect 15059 10724 15071 10727
rect 16132 10724 16160 10755
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18693 10795 18751 10801
rect 18693 10792 18705 10795
rect 18104 10764 18705 10792
rect 18104 10752 18110 10764
rect 18693 10761 18705 10764
rect 18739 10761 18751 10795
rect 18693 10755 18751 10761
rect 17221 10727 17279 10733
rect 17221 10724 17233 10727
rect 15059 10696 15792 10724
rect 16132 10696 17233 10724
rect 15059 10693 15071 10696
rect 15013 10687 15071 10693
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 5813 10619 5871 10625
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10588 4951 10591
rect 5442 10588 5448 10600
rect 4939 10560 5448 10588
rect 4939 10557 4951 10560
rect 4893 10551 4951 10557
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5828 10588 5856 10619
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 11698 10656 11704 10668
rect 11659 10628 11704 10656
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 15194 10656 15200 10668
rect 15151 10628 15200 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 8202 10588 8208 10600
rect 5828 10560 8208 10588
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8570 10588 8576 10600
rect 8531 10560 8576 10588
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 9398 10588 9404 10600
rect 9359 10560 9404 10588
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 10744 10560 11897 10588
rect 10744 10548 10750 10560
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 11885 10551 11943 10557
rect 14384 10560 14473 10588
rect 9677 10523 9735 10529
rect 9677 10489 9689 10523
rect 9723 10520 9735 10523
rect 12618 10520 12624 10532
rect 9723 10492 12624 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2924 10424 2973 10452
rect 2924 10412 2930 10424
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4525 10455 4583 10461
rect 4525 10452 4537 10455
rect 4488 10424 4537 10452
rect 4488 10412 4494 10424
rect 4525 10421 4537 10424
rect 4571 10421 4583 10455
rect 10870 10452 10876 10464
rect 10831 10424 10876 10452
rect 4525 10415 4583 10421
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 14384 10452 14412 10560
rect 14461 10557 14473 10560
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 14936 10520 14964 10619
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15764 10665 15792 10696
rect 17221 10693 17233 10696
rect 17267 10693 17279 10727
rect 17221 10687 17279 10693
rect 17954 10684 17960 10736
rect 18012 10684 18018 10736
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 15378 10548 15384 10600
rect 15436 10588 15442 10600
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 15436 10560 15669 10588
rect 15436 10548 15442 10560
rect 15657 10557 15669 10560
rect 15703 10557 15715 10591
rect 15657 10551 15715 10557
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16850 10588 16856 10600
rect 16632 10560 16856 10588
rect 16632 10548 16638 10560
rect 16850 10548 16856 10560
rect 16908 10588 16914 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16908 10560 16957 10588
rect 16908 10548 16914 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 17218 10588 17224 10600
rect 16945 10551 17003 10557
rect 17052 10560 17224 10588
rect 15470 10520 15476 10532
rect 14936 10492 15476 10520
rect 15470 10480 15476 10492
rect 15528 10520 15534 10532
rect 17052 10520 17080 10560
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 15528 10492 17080 10520
rect 15528 10480 15534 10492
rect 14148 10424 14412 10452
rect 14148 10412 14154 10424
rect 1104 10362 19412 10384
rect 1104 10310 4001 10362
rect 4053 10310 4065 10362
rect 4117 10310 4129 10362
rect 4181 10310 4193 10362
rect 4245 10310 4257 10362
rect 4309 10310 10104 10362
rect 10156 10310 10168 10362
rect 10220 10310 10232 10362
rect 10284 10310 10296 10362
rect 10348 10310 10360 10362
rect 10412 10310 16206 10362
rect 16258 10310 16270 10362
rect 16322 10310 16334 10362
rect 16386 10310 16398 10362
rect 16450 10310 16462 10362
rect 16514 10310 19412 10362
rect 1104 10288 19412 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2774 10248 2780 10260
rect 1903 10220 2780 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5537 10251 5595 10257
rect 5537 10248 5549 10251
rect 5500 10220 5549 10248
rect 5500 10208 5506 10220
rect 5537 10217 5549 10220
rect 5583 10217 5595 10251
rect 10686 10248 10692 10260
rect 10647 10220 10692 10248
rect 5537 10211 5595 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 11406 10251 11464 10257
rect 11406 10248 11418 10251
rect 10928 10220 11418 10248
rect 10928 10208 10934 10220
rect 11406 10217 11418 10220
rect 11452 10217 11464 10251
rect 11406 10211 11464 10217
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18049 10251 18107 10257
rect 18049 10248 18061 10251
rect 18012 10220 18061 10248
rect 18012 10208 18018 10220
rect 18049 10217 18061 10220
rect 18095 10217 18107 10251
rect 18049 10211 18107 10217
rect 3786 10180 3792 10192
rect 2976 10152 3792 10180
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2976 10121 3004 10152
rect 3786 10140 3792 10152
rect 3844 10140 3850 10192
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10081 3019 10115
rect 6914 10112 6920 10124
rect 6875 10084 6920 10112
rect 2961 10075 3019 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 8386 10112 8392 10124
rect 7147 10084 8392 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 8570 10072 8576 10124
rect 8628 10112 8634 10124
rect 8938 10112 8944 10124
rect 8628 10084 8944 10112
rect 8628 10072 8634 10084
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 12894 10112 12900 10124
rect 11195 10084 12900 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 15378 10112 15384 10124
rect 15339 10084 15384 10112
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15528 10084 15573 10112
rect 15528 10072 15534 10084
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3752 10016 3801 10044
rect 3752 10004 3758 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 7009 10047 7067 10053
rect 7009 10044 7021 10047
rect 6052 10016 7021 10044
rect 6052 10004 6058 10016
rect 7009 10013 7021 10016
rect 7055 10013 7067 10047
rect 7009 10007 7067 10013
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7374 10044 7380 10056
rect 7239 10016 7380 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 15565 10047 15623 10053
rect 15565 10044 15577 10047
rect 14783 10016 15577 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 15565 10013 15577 10016
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 4062 9976 4068 9988
rect 4023 9948 4068 9976
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 4522 9936 4528 9988
rect 4580 9936 4586 9988
rect 6181 9979 6239 9985
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 7834 9976 7840 9988
rect 6227 9948 7840 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 7834 9936 7840 9948
rect 7892 9936 7898 9988
rect 9214 9976 9220 9988
rect 9175 9948 9220 9976
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9950 9936 9956 9988
rect 10008 9936 10014 9988
rect 12434 9936 12440 9988
rect 12492 9936 12498 9988
rect 13998 9936 14004 9988
rect 14056 9976 14062 9988
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 14056 9948 14565 9976
rect 14056 9936 14062 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 15580 9976 15608 10007
rect 15654 10004 15660 10056
rect 15712 10044 15718 10056
rect 15712 10016 15757 10044
rect 15712 10004 15718 10016
rect 16758 10004 16764 10056
rect 16816 10044 16822 10056
rect 17313 10047 17371 10053
rect 17313 10044 17325 10047
rect 16816 10016 17325 10044
rect 16816 10004 16822 10016
rect 17313 10013 17325 10016
rect 17359 10044 17371 10047
rect 17957 10047 18015 10053
rect 17957 10044 17969 10047
rect 17359 10016 17969 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 17957 10013 17969 10016
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 16022 9976 16028 9988
rect 15580 9948 16028 9976
rect 14553 9939 14611 9945
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 6086 9908 6092 9920
rect 6047 9880 6092 9908
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 6730 9908 6736 9920
rect 6691 9880 6736 9908
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 12897 9911 12955 9917
rect 12897 9908 12909 9911
rect 11756 9880 12909 9908
rect 11756 9868 11762 9880
rect 12897 9877 12909 9880
rect 12943 9877 12955 9911
rect 12897 9871 12955 9877
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15197 9911 15255 9917
rect 15197 9908 15209 9911
rect 14976 9880 15209 9908
rect 14976 9868 14982 9880
rect 15197 9877 15209 9880
rect 15243 9877 15255 9911
rect 15197 9871 15255 9877
rect 17405 9911 17463 9917
rect 17405 9877 17417 9911
rect 17451 9908 17463 9911
rect 18138 9908 18144 9920
rect 17451 9880 18144 9908
rect 17451 9877 17463 9880
rect 17405 9871 17463 9877
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 1104 9818 19412 9840
rect 1104 9766 7052 9818
rect 7104 9766 7116 9818
rect 7168 9766 7180 9818
rect 7232 9766 7244 9818
rect 7296 9766 7308 9818
rect 7360 9766 13155 9818
rect 13207 9766 13219 9818
rect 13271 9766 13283 9818
rect 13335 9766 13347 9818
rect 13399 9766 13411 9818
rect 13463 9766 19412 9818
rect 1104 9744 19412 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 1765 9707 1823 9713
rect 1765 9704 1777 9707
rect 1636 9676 1777 9704
rect 1636 9664 1642 9676
rect 1765 9673 1777 9676
rect 1811 9673 1823 9707
rect 1765 9667 1823 9673
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 3881 9707 3939 9713
rect 3752 9676 3832 9704
rect 3752 9664 3758 9676
rect 3804 9636 3832 9676
rect 3881 9673 3893 9707
rect 3927 9704 3939 9707
rect 4062 9704 4068 9716
rect 3927 9676 4068 9704
rect 3927 9673 3939 9676
rect 3881 9667 3939 9673
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 9214 9704 9220 9716
rect 9175 9676 9220 9704
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 15654 9704 15660 9716
rect 15615 9676 15660 9704
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 6641 9639 6699 9645
rect 3252 9608 3740 9636
rect 3804 9608 6408 9636
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1544 9540 1685 9568
rect 1544 9528 1550 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 2130 9568 2136 9580
rect 1903 9540 2136 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 2130 9528 2136 9540
rect 2188 9568 2194 9580
rect 2958 9568 2964 9580
rect 2188 9540 2964 9568
rect 2188 9528 2194 9540
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 3252 9500 3280 9608
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3384 9540 3617 9568
rect 3384 9528 3390 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3712 9568 3740 9608
rect 4430 9568 4436 9580
rect 3712 9540 4436 9568
rect 3605 9531 3663 9537
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 5442 9568 5448 9580
rect 4755 9540 5448 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 6380 9577 6408 9608
rect 6641 9605 6653 9639
rect 6687 9636 6699 9639
rect 6730 9636 6736 9648
rect 6687 9608 6736 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 6730 9596 6736 9608
rect 6788 9596 6794 9648
rect 7190 9596 7196 9648
rect 7248 9596 7254 9648
rect 9582 9636 9588 9648
rect 9508 9608 9588 9636
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 9398 9568 9404 9580
rect 9359 9540 9404 9568
rect 6365 9531 6423 9537
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 9508 9577 9536 9608
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 10686 9596 10692 9648
rect 10744 9596 10750 9648
rect 13998 9636 14004 9648
rect 12820 9608 14004 9636
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 10704 9568 10732 9596
rect 12820 9577 12848 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 14734 9596 14740 9648
rect 14792 9596 14798 9648
rect 18138 9596 18144 9648
rect 18196 9596 18202 9648
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10704 9540 10793 9568
rect 9493 9531 9551 9537
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9537 12863 9571
rect 15838 9568 15844 9580
rect 15799 9540 15844 9568
rect 12805 9531 12863 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3252 9472 3433 9500
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9500 3755 9503
rect 3786 9500 3792 9512
rect 3743 9472 3792 9500
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 3528 9364 3556 9463
rect 3786 9460 3792 9472
rect 3844 9500 3850 9512
rect 4341 9503 4399 9509
rect 4341 9500 4353 9503
rect 3844 9472 4353 9500
rect 3844 9460 3850 9472
rect 4341 9469 4353 9472
rect 4387 9469 4399 9503
rect 4798 9500 4804 9512
rect 4759 9472 4804 9500
rect 4341 9463 4399 9469
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 9030 9500 9036 9512
rect 8444 9472 9036 9500
rect 8444 9460 8450 9472
rect 9030 9460 9036 9472
rect 9088 9500 9094 9512
rect 9585 9503 9643 9509
rect 9585 9500 9597 9503
rect 9088 9472 9597 9500
rect 9088 9460 9094 9472
rect 9585 9469 9597 9472
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9500 10931 9503
rect 11698 9500 11704 9512
rect 10919 9472 11704 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 9692 9432 9720 9463
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9500 13507 9503
rect 13725 9503 13783 9509
rect 13495 9472 13584 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 11514 9432 11520 9444
rect 9692 9404 11520 9432
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 4338 9364 4344 9376
rect 2280 9336 4344 9364
rect 2280 9324 2286 9336
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 8110 9364 8116 9376
rect 8071 9336 8116 9364
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9456 9336 10425 9364
rect 9456 9324 9462 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 12621 9367 12679 9373
rect 12621 9364 12633 9367
rect 12584 9336 12633 9364
rect 12584 9324 12590 9336
rect 12621 9333 12633 9336
rect 12667 9333 12679 9367
rect 13556 9364 13584 9472
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 14918 9500 14924 9512
rect 13771 9472 14924 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15102 9460 15108 9512
rect 15160 9500 15166 9512
rect 15197 9503 15255 9509
rect 15197 9500 15209 9503
rect 15160 9472 15209 9500
rect 15160 9460 15166 9472
rect 15197 9469 15209 9472
rect 15243 9500 15255 9503
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15243 9472 16037 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 16850 9500 16856 9512
rect 16811 9472 16856 9500
rect 16025 9463 16083 9469
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 17126 9500 17132 9512
rect 17087 9472 17132 9500
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 14090 9364 14096 9376
rect 13556 9336 14096 9364
rect 12621 9327 12679 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 18506 9324 18512 9376
rect 18564 9364 18570 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 18564 9336 18613 9364
rect 18564 9324 18570 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18601 9327 18659 9333
rect 1104 9274 19412 9296
rect 1104 9222 4001 9274
rect 4053 9222 4065 9274
rect 4117 9222 4129 9274
rect 4181 9222 4193 9274
rect 4245 9222 4257 9274
rect 4309 9222 10104 9274
rect 10156 9222 10168 9274
rect 10220 9222 10232 9274
rect 10284 9222 10296 9274
rect 10348 9222 10360 9274
rect 10412 9222 16206 9274
rect 16258 9222 16270 9274
rect 16322 9222 16334 9274
rect 16386 9222 16398 9274
rect 16450 9222 16462 9274
rect 16514 9222 19412 9274
rect 1104 9200 19412 9222
rect 4157 9163 4215 9169
rect 4157 9129 4169 9163
rect 4203 9160 4215 9163
rect 4522 9160 4528 9172
rect 4203 9132 4528 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7101 9163 7159 9169
rect 7101 9160 7113 9163
rect 6972 9132 7113 9160
rect 6972 9120 6978 9132
rect 7101 9129 7113 9132
rect 7147 9129 7159 9163
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 7101 9123 7159 9129
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 12406 9132 13185 9160
rect 6549 9095 6607 9101
rect 6549 9061 6561 9095
rect 6595 9092 6607 9095
rect 7190 9092 7196 9104
rect 6595 9064 7196 9092
rect 6595 9061 6607 9064
rect 6549 9055 6607 9061
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 8294 9024 8300 9036
rect 7607 8996 8300 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 5258 8956 5264 8968
rect 4111 8928 5264 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 5258 8916 5264 8928
rect 5316 8956 5322 8968
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 5316 8928 5641 8956
rect 5316 8916 5322 8928
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 6454 8956 6460 8968
rect 6415 8928 6460 8956
rect 5629 8919 5687 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 8110 8956 8116 8968
rect 7515 8928 8116 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 11054 8956 11060 8968
rect 10091 8928 11060 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8956 12127 8959
rect 12406 8956 12434 9132
rect 13173 9129 13185 9132
rect 13219 9160 13231 9163
rect 14826 9160 14832 9172
rect 13219 9132 14832 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 14826 9120 14832 9132
rect 14884 9120 14890 9172
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 15473 9163 15531 9169
rect 15473 9160 15485 9163
rect 15436 9132 15485 9160
rect 15436 9120 15442 9132
rect 15473 9129 15485 9132
rect 15519 9129 15531 9163
rect 15473 9123 15531 9129
rect 16945 9163 17003 9169
rect 16945 9129 16957 9163
rect 16991 9160 17003 9163
rect 17126 9160 17132 9172
rect 16991 9132 17132 9160
rect 16991 9129 17003 9132
rect 16945 9123 17003 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 15838 9092 15844 9104
rect 15212 9064 15844 9092
rect 15212 9033 15240 9064
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 15197 9027 15255 9033
rect 15197 8993 15209 9027
rect 15243 8993 15255 9027
rect 15197 8987 15255 8993
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 17221 9027 17279 9033
rect 17221 9024 17233 9027
rect 16632 8996 17233 9024
rect 16632 8984 16638 8996
rect 17221 8993 17233 8996
rect 17267 9024 17279 9027
rect 17586 9024 17592 9036
rect 17267 8996 17592 9024
rect 17267 8993 17279 8996
rect 17221 8987 17279 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 18506 9024 18512 9036
rect 18467 8996 18512 9024
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 14182 8956 14188 8968
rect 12115 8928 12434 8956
rect 14143 8928 14188 8956
rect 12115 8925 12127 8928
rect 12069 8919 12127 8925
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 15102 8956 15108 8968
rect 15063 8928 15108 8956
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15620 8928 16129 8956
rect 15620 8916 15626 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 17126 8956 17132 8968
rect 17087 8928 17132 8956
rect 16117 8919 16175 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8956 17463 8959
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 17451 8928 18153 8956
rect 17451 8925 17463 8928
rect 17405 8919 17463 8925
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8956 18383 8959
rect 18690 8956 18696 8968
rect 18371 8928 18696 8956
rect 18371 8925 18383 8928
rect 18325 8919 18383 8925
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 4709 8891 4767 8897
rect 4709 8888 4721 8891
rect 3752 8860 4721 8888
rect 3752 8848 3758 8860
rect 4709 8857 4721 8860
rect 4755 8857 4767 8891
rect 4709 8851 4767 8857
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8888 4951 8891
rect 6086 8888 6092 8900
rect 4939 8860 6092 8888
rect 4939 8857 4951 8860
rect 4893 8851 4951 8857
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8888 13323 8891
rect 13814 8888 13820 8900
rect 13311 8860 13820 8888
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 16022 8848 16028 8900
rect 16080 8888 16086 8900
rect 17328 8888 17356 8919
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 16080 8860 17356 8888
rect 16080 8848 16086 8860
rect 5534 8820 5540 8832
rect 5495 8792 5540 8820
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11112 8792 11897 8820
rect 11112 8780 11118 8792
rect 11885 8789 11897 8792
rect 11931 8820 11943 8823
rect 12342 8820 12348 8832
rect 11931 8792 12348 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 14274 8820 14280 8832
rect 14235 8792 14280 8820
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 14424 8792 15945 8820
rect 14424 8780 14430 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 15933 8783 15991 8789
rect 1104 8730 19412 8752
rect 1104 8678 7052 8730
rect 7104 8678 7116 8730
rect 7168 8678 7180 8730
rect 7232 8678 7244 8730
rect 7296 8678 7308 8730
rect 7360 8678 13155 8730
rect 13207 8678 13219 8730
rect 13271 8678 13283 8730
rect 13335 8678 13347 8730
rect 13399 8678 13411 8730
rect 13463 8678 19412 8730
rect 1104 8656 19412 8678
rect 6454 8576 6460 8628
rect 6512 8616 6518 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6512 8588 6561 8616
rect 6512 8576 6518 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 6549 8579 6607 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 14366 8616 14372 8628
rect 7616 8588 8432 8616
rect 7616 8576 7622 8588
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3292 8520 3985 8548
rect 3292 8508 3298 8520
rect 3973 8517 3985 8520
rect 4019 8517 4031 8551
rect 5534 8548 5540 8560
rect 5198 8520 5540 8548
rect 3973 8511 4031 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 2038 8480 2044 8492
rect 1728 8452 2044 8480
rect 1728 8440 1734 8452
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 2222 8440 2228 8452
rect 2280 8480 2286 8492
rect 2682 8480 2688 8492
rect 2280 8452 2688 8480
rect 2280 8440 2286 8452
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 1486 8372 1492 8424
rect 1544 8412 1550 8424
rect 2133 8415 2191 8421
rect 2133 8412 2145 8415
rect 1544 8384 2145 8412
rect 1544 8372 1550 8384
rect 2133 8381 2145 8384
rect 2179 8381 2191 8415
rect 2133 8375 2191 8381
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 2869 8415 2927 8421
rect 2869 8412 2881 8415
rect 2363 8384 2881 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 2869 8381 2881 8384
rect 2915 8381 2927 8415
rect 3068 8412 3096 8443
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3200 8452 3245 8480
rect 3200 8440 3206 8452
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6236 8452 6377 8480
rect 6236 8440 6242 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 8110 8480 8116 8492
rect 7791 8452 8116 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 3234 8412 3240 8424
rect 3068 8384 3240 8412
rect 2869 8375 2927 8381
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 3694 8412 3700 8424
rect 3655 8384 3700 8412
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 5442 8344 5448 8356
rect 5403 8316 5448 8344
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 6380 8344 6408 8443
rect 7576 8412 7604 8443
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8404 8489 8432 8588
rect 13280 8588 14372 8616
rect 12802 8508 12808 8560
rect 12860 8508 12866 8560
rect 13280 8557 13308 8588
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 15436 8588 16681 8616
rect 15436 8576 15442 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 13265 8551 13323 8557
rect 13265 8517 13277 8551
rect 13311 8517 13323 8551
rect 13265 8511 13323 8517
rect 14185 8551 14243 8557
rect 14185 8517 14197 8551
rect 14231 8548 14243 8551
rect 14274 8548 14280 8560
rect 14231 8520 14280 8548
rect 14231 8517 14243 8520
rect 14185 8511 14243 8517
rect 14274 8508 14280 8520
rect 14332 8548 14338 8560
rect 14829 8551 14887 8557
rect 14829 8548 14841 8551
rect 14332 8520 14841 8548
rect 14332 8508 14338 8520
rect 14829 8517 14841 8520
rect 14875 8517 14887 8551
rect 14829 8511 14887 8517
rect 16025 8551 16083 8557
rect 16025 8517 16037 8551
rect 16071 8548 16083 8551
rect 16071 8520 17080 8548
rect 16071 8517 16083 8520
rect 16025 8511 16083 8517
rect 8389 8483 8447 8489
rect 8260 8452 8305 8480
rect 8260 8440 8266 8452
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 8662 8480 8668 8492
rect 8435 8452 8668 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11054 8480 11060 8492
rect 10827 8452 11060 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15252 8452 15945 8480
rect 15252 8440 15258 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8480 16175 8483
rect 16574 8480 16580 8492
rect 16163 8452 16580 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 17052 8489 17080 8520
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 18506 8480 18512 8492
rect 18371 8452 18512 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 8294 8412 8300 8424
rect 7576 8384 8300 8412
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 12710 8412 12716 8424
rect 11839 8384 12716 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 17126 8412 17132 8424
rect 17039 8384 17132 8412
rect 13541 8375 13599 8381
rect 9950 8344 9956 8356
rect 6380 8316 9956 8344
rect 9950 8304 9956 8316
rect 10008 8304 10014 8356
rect 10873 8347 10931 8353
rect 10873 8313 10885 8347
rect 10919 8344 10931 8347
rect 11238 8344 11244 8356
rect 10919 8316 11244 8344
rect 10919 8313 10931 8316
rect 10873 8307 10931 8313
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 13556 8344 13584 8375
rect 17126 8372 17132 8384
rect 17184 8412 17190 8424
rect 17957 8415 18015 8421
rect 17957 8412 17969 8415
rect 17184 8384 17969 8412
rect 17184 8372 17190 8384
rect 17957 8381 17969 8384
rect 18003 8381 18015 8415
rect 17957 8375 18015 8381
rect 18417 8415 18475 8421
rect 18417 8381 18429 8415
rect 18463 8412 18475 8415
rect 18690 8412 18696 8424
rect 18463 8384 18696 8412
rect 18463 8381 18475 8384
rect 18417 8375 18475 8381
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 13722 8344 13728 8356
rect 13556 8316 13728 8344
rect 1670 8236 1676 8288
rect 1728 8276 1734 8288
rect 1857 8279 1915 8285
rect 1857 8276 1869 8279
rect 1728 8248 1869 8276
rect 1728 8236 1734 8248
rect 1857 8245 1869 8248
rect 1903 8245 1915 8279
rect 1857 8239 1915 8245
rect 8297 8279 8355 8285
rect 8297 8245 8309 8279
rect 8343 8276 8355 8279
rect 8754 8276 8760 8288
rect 8343 8248 8760 8276
rect 8343 8245 8355 8248
rect 8297 8239 8355 8245
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13556 8276 13584 8316
rect 13722 8304 13728 8316
rect 13780 8344 13786 8356
rect 14001 8347 14059 8353
rect 14001 8344 14013 8347
rect 13780 8316 14013 8344
rect 13780 8304 13786 8316
rect 14001 8313 14013 8316
rect 14047 8313 14059 8347
rect 14001 8307 14059 8313
rect 14090 8304 14096 8356
rect 14148 8344 14154 8356
rect 15013 8347 15071 8353
rect 15013 8344 15025 8347
rect 14148 8316 15025 8344
rect 14148 8304 14154 8316
rect 15013 8313 15025 8316
rect 15059 8344 15071 8347
rect 15059 8316 16988 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 16960 8288 16988 8316
rect 12952 8248 13584 8276
rect 12952 8236 12958 8248
rect 16942 8236 16948 8288
rect 17000 8236 17006 8288
rect 1104 8186 19412 8208
rect 1104 8134 4001 8186
rect 4053 8134 4065 8186
rect 4117 8134 4129 8186
rect 4181 8134 4193 8186
rect 4245 8134 4257 8186
rect 4309 8134 10104 8186
rect 10156 8134 10168 8186
rect 10220 8134 10232 8186
rect 10284 8134 10296 8186
rect 10348 8134 10360 8186
rect 10412 8134 16206 8186
rect 16258 8134 16270 8186
rect 16322 8134 16334 8186
rect 16386 8134 16398 8186
rect 16450 8134 16462 8186
rect 16514 8134 19412 8186
rect 1104 8112 19412 8134
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6420 8044 6745 8072
rect 6420 8032 6426 8044
rect 6733 8041 6745 8044
rect 6779 8072 6791 8075
rect 6779 8044 7880 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 6454 8004 6460 8016
rect 5920 7976 6460 8004
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 5920 7877 5948 7976
rect 6454 7964 6460 7976
rect 6512 7964 6518 8016
rect 7852 8004 7880 8044
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 10689 8075 10747 8081
rect 10689 8072 10701 8075
rect 8352 8044 10701 8072
rect 8352 8032 8358 8044
rect 10689 8041 10701 8044
rect 10735 8041 10747 8075
rect 10689 8035 10747 8041
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 12860 8044 13461 8072
rect 12860 8032 12866 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 15838 8072 15844 8084
rect 15799 8044 15844 8072
rect 13449 8035 13507 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 7852 7976 8984 8004
rect 8956 7948 8984 7976
rect 7558 7936 7564 7948
rect 7519 7908 7564 7936
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7905 7711 7939
rect 8938 7936 8944 7948
rect 8899 7908 8944 7936
rect 7653 7899 7711 7905
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 3326 7800 3332 7812
rect 2898 7772 3332 7800
rect 3326 7760 3332 7772
rect 3384 7760 3390 7812
rect 4816 7800 4844 7831
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6144 7840 6653 7868
rect 6144 7828 6150 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 7432 7840 7481 7868
rect 7432 7828 7438 7840
rect 7469 7837 7481 7840
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 6178 7800 6184 7812
rect 4816 7772 6184 7800
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 3142 7732 3148 7744
rect 3103 7704 3148 7732
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5258 7732 5264 7744
rect 5031 7704 5264 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5994 7732 6000 7744
rect 5955 7704 6000 7732
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 6696 7704 7297 7732
rect 6696 7692 6702 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7668 7732 7696 7899
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 12618 7936 12624 7948
rect 12579 7908 12624 7936
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12894 7936 12900 7948
rect 12855 7908 12900 7936
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 14090 7936 14096 7948
rect 14051 7908 14096 7936
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7936 14427 7939
rect 15378 7936 15384 7948
rect 14415 7908 15384 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 7800 7840 7845 7868
rect 7800 7828 7806 7840
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 13357 7871 13415 7877
rect 13357 7868 13369 7871
rect 13044 7840 13369 7868
rect 13044 7828 13050 7840
rect 13357 7837 13369 7840
rect 13403 7837 13415 7871
rect 13357 7831 13415 7837
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 18196 7840 18245 7868
rect 18196 7828 18202 7840
rect 18233 7837 18245 7840
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 9122 7760 9128 7812
rect 9180 7800 9186 7812
rect 9217 7803 9275 7809
rect 9217 7800 9229 7803
rect 9180 7772 9229 7800
rect 9180 7760 9186 7772
rect 9217 7769 9229 7772
rect 9263 7769 9275 7803
rect 10594 7800 10600 7812
rect 10442 7772 10600 7800
rect 9217 7763 9275 7769
rect 10594 7760 10600 7772
rect 10652 7760 10658 7812
rect 11238 7760 11244 7812
rect 11296 7800 11302 7812
rect 11296 7772 11454 7800
rect 11296 7760 11302 7772
rect 9030 7732 9036 7744
rect 7668 7704 9036 7732
rect 7285 7695 7343 7701
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11149 7735 11207 7741
rect 11149 7732 11161 7735
rect 10928 7704 11161 7732
rect 10928 7692 10934 7704
rect 11149 7701 11161 7704
rect 11195 7701 11207 7735
rect 11149 7695 11207 7701
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18230 7732 18236 7744
rect 18187 7704 18236 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 1104 7642 19412 7664
rect 1104 7590 7052 7642
rect 7104 7590 7116 7642
rect 7168 7590 7180 7642
rect 7232 7590 7244 7642
rect 7296 7590 7308 7642
rect 7360 7590 13155 7642
rect 13207 7590 13219 7642
rect 13271 7590 13283 7642
rect 13335 7590 13347 7642
rect 13399 7590 13411 7642
rect 13463 7590 19412 7642
rect 1104 7568 19412 7590
rect 3326 7528 3332 7540
rect 3287 7500 3332 7528
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 9122 7528 9128 7540
rect 6052 7500 6960 7528
rect 9083 7500 9128 7528
rect 6052 7488 6058 7500
rect 6638 7460 6644 7472
rect 6599 7432 6644 7460
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 6932 7460 6960 7500
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 9950 7528 9956 7540
rect 9911 7500 9956 7528
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10594 7488 10600 7540
rect 10652 7528 10658 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 10652 7500 10701 7528
rect 10652 7488 10658 7500
rect 10689 7497 10701 7500
rect 10735 7497 10747 7531
rect 10689 7491 10747 7497
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 14829 7531 14887 7537
rect 14829 7528 14841 7531
rect 14792 7500 14841 7528
rect 14792 7488 14798 7500
rect 14829 7497 14841 7500
rect 14875 7497 14887 7531
rect 15470 7528 15476 7540
rect 15431 7500 15476 7528
rect 14829 7491 14887 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 18138 7528 18144 7540
rect 15580 7500 18144 7528
rect 6932 7432 7130 7460
rect 9582 7420 9588 7472
rect 9640 7460 9646 7472
rect 9640 7432 10824 7460
rect 9640 7420 9646 7432
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 3142 7392 3148 7404
rect 2639 7364 3148 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7361 3479 7395
rect 8754 7392 8760 7404
rect 8715 7364 8760 7392
rect 3421 7355 3479 7361
rect 2038 7284 2044 7336
rect 2096 7324 2102 7336
rect 2225 7327 2283 7333
rect 2225 7324 2237 7327
rect 2096 7296 2237 7324
rect 2096 7284 2102 7296
rect 2225 7293 2237 7296
rect 2271 7293 2283 7327
rect 2225 7287 2283 7293
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 3234 7324 3240 7336
rect 2731 7296 3240 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 3436 7200 3464 7355
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 10796 7401 10824 7432
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 6362 7324 6368 7336
rect 6323 7296 6368 7324
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 7432 7296 8677 7324
rect 7432 7284 7438 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 10060 7324 10088 7355
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12768 7364 13001 7392
rect 12768 7352 12774 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13814 7392 13820 7404
rect 13136 7364 13181 7392
rect 13727 7364 13820 7392
rect 13136 7352 13142 7364
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 10962 7324 10968 7336
rect 10060 7296 10968 7324
rect 8665 7287 8723 7293
rect 10962 7284 10968 7296
rect 11020 7324 11026 7336
rect 13832 7324 13860 7352
rect 11020 7296 13860 7324
rect 14936 7324 14964 7355
rect 15010 7352 15016 7404
rect 15068 7392 15074 7404
rect 15580 7401 15608 7500
rect 18138 7488 18144 7500
rect 18196 7488 18202 7540
rect 18690 7528 18696 7540
rect 18651 7500 18696 7528
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 18230 7420 18236 7472
rect 18288 7420 18294 7472
rect 15565 7395 15623 7401
rect 15565 7392 15577 7395
rect 15068 7364 15577 7392
rect 15068 7352 15074 7364
rect 15565 7361 15577 7364
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 16758 7324 16764 7336
rect 14936 7296 16764 7324
rect 11020 7284 11026 7296
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 16942 7324 16948 7336
rect 16903 7296 16948 7324
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 17218 7324 17224 7336
rect 17179 7296 17224 7324
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 12986 7256 12992 7268
rect 7668 7228 12434 7256
rect 3418 7188 3424 7200
rect 3331 7160 3424 7188
rect 3418 7148 3424 7160
rect 3476 7188 3482 7200
rect 7668 7188 7696 7228
rect 8110 7188 8116 7200
rect 3476 7160 7696 7188
rect 8071 7160 8116 7188
rect 3476 7148 3482 7160
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 12406 7188 12434 7228
rect 12636 7228 12992 7256
rect 12636 7188 12664 7228
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 12802 7188 12808 7200
rect 12406 7160 12664 7188
rect 12763 7160 12808 7188
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 14001 7191 14059 7197
rect 14001 7157 14013 7191
rect 14047 7188 14059 7191
rect 15010 7188 15016 7200
rect 14047 7160 15016 7188
rect 14047 7157 14059 7160
rect 14001 7151 14059 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 1104 7098 19412 7120
rect 1104 7046 4001 7098
rect 4053 7046 4065 7098
rect 4117 7046 4129 7098
rect 4181 7046 4193 7098
rect 4245 7046 4257 7098
rect 4309 7046 10104 7098
rect 10156 7046 10168 7098
rect 10220 7046 10232 7098
rect 10284 7046 10296 7098
rect 10348 7046 10360 7098
rect 10412 7046 16206 7098
rect 16258 7046 16270 7098
rect 16322 7046 16334 7098
rect 16386 7046 16398 7098
rect 16450 7046 16462 7098
rect 16514 7046 19412 7098
rect 1104 7024 19412 7046
rect 7374 6984 7380 6996
rect 7335 6956 7380 6984
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 9582 6984 9588 6996
rect 9543 6956 9588 6984
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 16114 6916 16120 6928
rect 15948 6888 16120 6916
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 3694 6848 3700 6860
rect 1452 6820 3700 6848
rect 1452 6808 1458 6820
rect 3694 6808 3700 6820
rect 3752 6848 3758 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3752 6820 3801 6848
rect 3752 6808 3758 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 7834 6848 7840 6860
rect 7795 6820 7840 6848
rect 3789 6811 3847 6817
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12710 6848 12716 6860
rect 12492 6820 12537 6848
rect 12671 6820 12716 6848
rect 12492 6808 12498 6820
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6848 15899 6851
rect 15948 6848 15976 6888
rect 16114 6876 16120 6888
rect 16172 6916 16178 6928
rect 17218 6916 17224 6928
rect 16172 6888 16804 6916
rect 17179 6888 17224 6916
rect 16172 6876 16178 6888
rect 15887 6820 15976 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16776 6857 16804 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 16761 6851 16819 6857
rect 16080 6820 16125 6848
rect 16080 6808 16086 6820
rect 16761 6817 16773 6851
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8110 6780 8116 6792
rect 7791 6752 8116 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 9950 6780 9956 6792
rect 9815 6752 9956 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6780 12863 6783
rect 13078 6780 13084 6792
rect 12851 6752 13084 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 15010 6780 15016 6792
rect 14875 6752 15016 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15934 6783 15992 6789
rect 15934 6749 15946 6783
rect 15980 6749 15992 6783
rect 15934 6743 15992 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16666 6780 16672 6792
rect 16163 6752 16672 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 4062 6712 4068 6724
rect 4023 6684 4068 6712
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 6454 6712 6460 6724
rect 5290 6684 6460 6712
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 5534 6644 5540 6656
rect 5495 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 14918 6644 14924 6656
rect 14879 6616 14924 6644
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 15654 6644 15660 6656
rect 15615 6616 15660 6644
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 15948 6644 15976 6743
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 16868 6712 16896 6743
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 17678 6780 17684 6792
rect 17368 6752 17684 6780
rect 17368 6740 17374 6752
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6780 17923 6783
rect 18322 6780 18328 6792
rect 17911 6752 18328 6780
rect 17911 6749 17923 6752
rect 17865 6743 17923 6749
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 16868 6684 17785 6712
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17773 6675 17831 6681
rect 17880 6644 17908 6743
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 15948 6616 17908 6644
rect 1104 6554 19412 6576
rect 1104 6502 7052 6554
rect 7104 6502 7116 6554
rect 7168 6502 7180 6554
rect 7232 6502 7244 6554
rect 7296 6502 7308 6554
rect 7360 6502 13155 6554
rect 13207 6502 13219 6554
rect 13271 6502 13283 6554
rect 13335 6502 13347 6554
rect 13399 6502 13411 6554
rect 13463 6502 19412 6554
rect 1104 6480 19412 6502
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 4062 6440 4068 6452
rect 3927 6412 4068 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4338 6440 4344 6452
rect 4212 6412 4344 6440
rect 4212 6400 4218 6412
rect 4338 6400 4344 6412
rect 4396 6440 4402 6452
rect 4890 6440 4896 6452
rect 4396 6412 4896 6440
rect 4396 6400 4402 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 6454 6440 6460 6452
rect 6415 6412 6460 6440
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 7653 6443 7711 6449
rect 7653 6409 7665 6443
rect 7699 6440 7711 6443
rect 7742 6440 7748 6452
rect 7699 6412 7748 6440
rect 7699 6409 7711 6412
rect 7653 6403 7711 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 13136 6412 13277 6440
rect 13136 6400 13142 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 15654 6440 15660 6452
rect 13265 6403 13323 6409
rect 14200 6412 15660 6440
rect 2682 6332 2688 6384
rect 2740 6372 2746 6384
rect 14200 6381 14228 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 16666 6440 16672 6452
rect 16627 6412 16672 6440
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 14185 6375 14243 6381
rect 2740 6344 4292 6372
rect 2740 6332 2746 6344
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2130 6304 2136 6316
rect 1903 6276 2136 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 4154 6304 4160 6316
rect 4115 6276 4160 6304
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4264 6313 4292 6344
rect 14185 6341 14197 6375
rect 14231 6341 14243 6375
rect 14185 6335 14243 6341
rect 14918 6332 14924 6384
rect 14976 6332 14982 6384
rect 15746 6332 15752 6384
rect 15804 6372 15810 6384
rect 15804 6344 17540 6372
rect 15804 6332 15810 6344
rect 17512 6316 17540 6344
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5534 6304 5540 6316
rect 5307 6276 5540 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 7834 6304 7840 6316
rect 7795 6276 7840 6304
rect 6365 6267 6423 6273
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 5074 6236 5080 6248
rect 4387 6208 5080 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 4080 6168 4108 6199
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6236 5411 6239
rect 5442 6236 5448 6248
rect 5399 6208 5448 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 4430 6168 4436 6180
rect 4080 6140 4436 6168
rect 4430 6128 4436 6140
rect 4488 6168 4494 6180
rect 4893 6171 4951 6177
rect 4893 6168 4905 6171
rect 4488 6140 4905 6168
rect 4488 6128 4494 6140
rect 4893 6137 4905 6140
rect 4939 6137 4951 6171
rect 4893 6131 4951 6137
rect 5258 6128 5264 6180
rect 5316 6168 5322 6180
rect 6380 6168 6408 6267
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6304 8079 6307
rect 8110 6304 8116 6316
rect 8067 6276 8116 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 12894 6264 12900 6316
rect 12952 6264 12958 6316
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 13780 6276 13921 6304
rect 13780 6264 13786 6276
rect 13909 6273 13921 6276
rect 13955 6273 13967 6307
rect 16850 6304 16856 6316
rect 16811 6276 16856 6304
rect 13909 6267 13967 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17494 6304 17500 6316
rect 17407 6276 17500 6304
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 17678 6304 17684 6316
rect 17639 6276 17684 6304
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6205 11575 6239
rect 11517 6199 11575 6205
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 12342 6236 12348 6248
rect 11839 6208 12348 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 5316 6140 6408 6168
rect 5316 6128 5322 6140
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 1854 6100 1860 6112
rect 1811 6072 1860 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 11532 6100 11560 6199
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 13740 6168 13768 6264
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 15620 6208 15669 6236
rect 15620 6196 15626 6208
rect 15657 6205 15669 6208
rect 15703 6236 15715 6239
rect 17037 6239 17095 6245
rect 17037 6236 17049 6239
rect 15703 6208 17049 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 17037 6205 17049 6208
rect 17083 6205 17095 6239
rect 17037 6199 17095 6205
rect 13004 6140 13768 6168
rect 12526 6100 12532 6112
rect 11532 6072 12532 6100
rect 12526 6060 12532 6072
rect 12584 6100 12590 6112
rect 13004 6100 13032 6140
rect 12584 6072 13032 6100
rect 12584 6060 12590 6072
rect 17402 6060 17408 6112
rect 17460 6100 17466 6112
rect 17589 6103 17647 6109
rect 17589 6100 17601 6103
rect 17460 6072 17601 6100
rect 17460 6060 17466 6072
rect 17589 6069 17601 6072
rect 17635 6069 17647 6103
rect 17589 6063 17647 6069
rect 1104 6010 19412 6032
rect 1104 5958 4001 6010
rect 4053 5958 4065 6010
rect 4117 5958 4129 6010
rect 4181 5958 4193 6010
rect 4245 5958 4257 6010
rect 4309 5958 10104 6010
rect 10156 5958 10168 6010
rect 10220 5958 10232 6010
rect 10284 5958 10296 6010
rect 10348 5958 10360 6010
rect 10412 5958 16206 6010
rect 16258 5958 16270 6010
rect 16322 5958 16334 6010
rect 16386 5958 16398 6010
rect 16450 5958 16462 6010
rect 16514 5958 19412 6010
rect 1104 5936 19412 5958
rect 3234 5896 3240 5908
rect 3195 5868 3240 5896
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 5074 5896 5080 5908
rect 5035 5868 5080 5896
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 7892 5868 8309 5896
rect 7892 5856 7898 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 12342 5896 12348 5908
rect 12303 5868 12348 5896
rect 8297 5859 8355 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 15933 5899 15991 5905
rect 15933 5865 15945 5899
rect 15979 5896 15991 5899
rect 16114 5896 16120 5908
rect 15979 5868 16120 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 18693 5899 18751 5905
rect 18693 5896 18705 5899
rect 16908 5868 18705 5896
rect 16908 5856 16914 5868
rect 18693 5865 18705 5868
rect 18739 5865 18751 5899
rect 18693 5859 18751 5865
rect 12710 5828 12716 5840
rect 4080 5800 6684 5828
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 4080 5760 4108 5800
rect 2188 5732 4108 5760
rect 2188 5720 2194 5732
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 4080 5701 4108 5732
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5534 5760 5540 5772
rect 5491 5732 5540 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 6656 5760 6684 5800
rect 7852 5800 12716 5828
rect 7852 5760 7880 5800
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 6656 5732 7880 5760
rect 9306 5720 9312 5772
rect 9364 5760 9370 5772
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 9364 5732 9505 5760
rect 9364 5720 9370 5732
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12492 5732 12541 5760
rect 12492 5720 12498 5732
rect 12529 5729 12541 5732
rect 12575 5729 12587 5763
rect 12802 5760 12808 5772
rect 12763 5732 12808 5760
rect 12529 5723 12587 5729
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 16868 5760 16896 5856
rect 15703 5732 16896 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 1489 5695 1547 5701
rect 1489 5692 1501 5695
rect 1452 5664 1501 5692
rect 1452 5652 1458 5664
rect 1489 5661 1501 5664
rect 1535 5661 1547 5695
rect 1489 5655 1547 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4338 5692 4344 5704
rect 4295 5664 4344 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 6362 5652 6368 5704
rect 6420 5692 6426 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6420 5664 6561 5692
rect 6420 5652 6426 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 9398 5692 9404 5704
rect 9359 5664 9404 5692
rect 6549 5655 6607 5661
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 9585 5695 9643 5701
rect 9585 5661 9597 5695
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 9723 5664 10701 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10870 5692 10876 5704
rect 10831 5664 10876 5692
rect 10689 5655 10747 5661
rect 1762 5624 1768 5636
rect 1723 5596 1768 5624
rect 1762 5584 1768 5596
rect 1820 5584 1826 5636
rect 3510 5624 3516 5636
rect 2990 5596 3516 5624
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 6825 5627 6883 5633
rect 6825 5593 6837 5627
rect 6871 5624 6883 5627
rect 6914 5624 6920 5636
rect 6871 5596 6920 5624
rect 6871 5593 6883 5596
rect 6825 5587 6883 5593
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 7558 5584 7564 5636
rect 7616 5584 7622 5636
rect 9122 5584 9128 5636
rect 9180 5624 9186 5636
rect 9600 5624 9628 5655
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11054 5692 11060 5704
rect 11015 5664 11060 5692
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 9180 5596 9628 5624
rect 12636 5624 12664 5655
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 15562 5692 15568 5704
rect 12768 5664 12813 5692
rect 15523 5664 15568 5692
rect 12768 5652 12774 5664
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 16574 5652 16580 5704
rect 16632 5692 16638 5704
rect 16942 5692 16948 5704
rect 16632 5664 16948 5692
rect 16632 5652 16638 5664
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 18322 5652 18328 5704
rect 18380 5652 18386 5704
rect 17218 5624 17224 5636
rect 12636 5596 13584 5624
rect 17179 5596 17224 5624
rect 9180 5584 9186 5596
rect 13556 5568 13584 5596
rect 17218 5584 17224 5596
rect 17276 5584 17282 5636
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 4246 5556 4252 5568
rect 4203 5528 4252 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 9217 5559 9275 5565
rect 9217 5525 9229 5559
rect 9263 5556 9275 5559
rect 9398 5556 9404 5568
rect 9263 5528 9404 5556
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 15930 5556 15936 5568
rect 13596 5528 15936 5556
rect 13596 5516 13602 5528
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 1104 5466 19412 5488
rect 1104 5414 7052 5466
rect 7104 5414 7116 5466
rect 7168 5414 7180 5466
rect 7232 5414 7244 5466
rect 7296 5414 7308 5466
rect 7360 5414 13155 5466
rect 13207 5414 13219 5466
rect 13271 5414 13283 5466
rect 13335 5414 13347 5466
rect 13399 5414 13411 5466
rect 13463 5414 19412 5466
rect 1104 5392 19412 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 1762 5352 1768 5364
rect 1535 5324 1768 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 3510 5352 3516 5364
rect 3471 5324 3516 5352
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 10873 5355 10931 5361
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 11054 5352 11060 5364
rect 10919 5324 11060 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 17037 5355 17095 5361
rect 17037 5321 17049 5355
rect 17083 5352 17095 5355
rect 17218 5352 17224 5364
rect 17083 5324 17224 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 18322 5352 18328 5364
rect 18283 5324 18328 5352
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 5258 5284 5264 5296
rect 3620 5256 5264 5284
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 3620 5225 3648 5256
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 9398 5284 9404 5296
rect 9359 5256 9404 5284
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 10626 5256 11621 5284
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 13265 5287 13323 5293
rect 13265 5284 13277 5287
rect 11609 5247 11667 5253
rect 12360 5256 13277 5284
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 4246 5216 4252 5228
rect 4207 5188 4252 5216
rect 3605 5179 3663 5185
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 1949 5151 2007 5157
rect 1949 5117 1961 5151
rect 1995 5148 2007 5151
rect 2130 5148 2136 5160
rect 1995 5120 2136 5148
rect 1995 5117 2007 5120
rect 1949 5111 2007 5117
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 4430 5148 4436 5160
rect 4387 5120 4436 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 6932 5148 6960 5179
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 7064 5188 7113 5216
rect 7064 5176 7070 5188
rect 7101 5185 7113 5188
rect 7147 5216 7159 5219
rect 7650 5216 7656 5228
rect 7147 5188 7656 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8294 5216 8300 5228
rect 8255 5188 8300 5216
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 12360 5225 12388 5256
rect 13265 5253 13277 5256
rect 13311 5253 13323 5287
rect 13265 5247 13323 5253
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8996 5188 9137 5216
rect 8996 5176 9002 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 13538 5216 13544 5228
rect 13403 5188 13544 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 8202 5148 8208 5160
rect 6932 5120 8208 5148
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5148 8447 5151
rect 9490 5148 9496 5160
rect 8435 5120 9496 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 11532 5148 11560 5179
rect 9824 5120 11560 5148
rect 12253 5151 12311 5157
rect 9824 5108 9830 5120
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12434 5148 12440 5160
rect 12299 5120 12440 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 13188 5148 13216 5179
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 14918 5216 14924 5228
rect 14879 5188 14924 5216
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 17402 5216 17408 5228
rect 17363 5188 17408 5216
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 18230 5216 18236 5228
rect 18191 5188 18236 5216
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 14274 5148 14280 5160
rect 13188 5120 14280 5148
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 14734 5148 14740 5160
rect 14695 5120 14740 5148
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 17310 5148 17316 5160
rect 17271 5120 17316 5148
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 4617 5083 4675 5089
rect 4617 5049 4629 5083
rect 4663 5080 4675 5083
rect 5534 5080 5540 5092
rect 4663 5052 5540 5080
rect 4663 5049 4675 5052
rect 4617 5043 4675 5049
rect 5534 5040 5540 5052
rect 5592 5040 5598 5092
rect 12710 5080 12716 5092
rect 12671 5052 12716 5080
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 7009 5015 7067 5021
rect 7009 5012 7021 5015
rect 6604 4984 7021 5012
rect 6604 4972 6610 4984
rect 7009 4981 7021 4984
rect 7055 4981 7067 5015
rect 7009 4975 7067 4981
rect 8573 5015 8631 5021
rect 8573 4981 8585 5015
rect 8619 5012 8631 5015
rect 9950 5012 9956 5024
rect 8619 4984 9956 5012
rect 8619 4981 8631 4984
rect 8573 4975 8631 4981
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 15105 5015 15163 5021
rect 15105 4981 15117 5015
rect 15151 5012 15163 5015
rect 15286 5012 15292 5024
rect 15151 4984 15292 5012
rect 15151 4981 15163 4984
rect 15105 4975 15163 4981
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 1104 4922 19412 4944
rect 1104 4870 4001 4922
rect 4053 4870 4065 4922
rect 4117 4870 4129 4922
rect 4181 4870 4193 4922
rect 4245 4870 4257 4922
rect 4309 4870 10104 4922
rect 10156 4870 10168 4922
rect 10220 4870 10232 4922
rect 10284 4870 10296 4922
rect 10348 4870 10360 4922
rect 10412 4870 16206 4922
rect 16258 4870 16270 4922
rect 16322 4870 16334 4922
rect 16386 4870 16398 4922
rect 16450 4870 16462 4922
rect 16514 4870 19412 4922
rect 1104 4848 19412 4870
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 7616 4780 7665 4808
rect 7616 4768 7622 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 8294 4808 8300 4820
rect 8255 4780 8300 4808
rect 7653 4771 7711 4777
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 9548 4780 10425 4808
rect 9548 4768 9554 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 10413 4771 10471 4777
rect 12621 4811 12679 4817
rect 12621 4777 12633 4811
rect 12667 4808 12679 4811
rect 12894 4808 12900 4820
rect 12667 4780 12900 4808
rect 12667 4777 12679 4780
rect 12621 4771 12679 4777
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 6914 4740 6920 4752
rect 6875 4712 6920 4740
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 17494 4700 17500 4752
rect 17552 4700 17558 4752
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 1728 4644 2237 4672
rect 1728 4632 1734 4644
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4672 2375 4675
rect 2682 4672 2688 4684
rect 2363 4644 2688 4672
rect 2363 4641 2375 4644
rect 2317 4635 2375 4641
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 6638 4672 6644 4684
rect 6599 4644 6644 4672
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 9582 4672 9588 4684
rect 7576 4644 9588 4672
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 5258 4604 5264 4616
rect 2464 4576 2509 4604
rect 5219 4576 5264 4604
rect 2464 4564 2470 4576
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 7576 4613 7604 4644
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 10870 4672 10876 4684
rect 10831 4644 10876 4672
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 15010 4672 15016 4684
rect 13964 4644 14504 4672
rect 14971 4644 15016 4672
rect 13964 4632 13970 4644
rect 14476 4616 14504 4644
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 17405 4675 17463 4681
rect 17405 4641 17417 4675
rect 17451 4672 17463 4675
rect 17512 4672 17540 4700
rect 17451 4644 17540 4672
rect 17451 4641 17463 4644
rect 17405 4635 17463 4641
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7524 4576 7573 4604
rect 7524 4564 7530 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 8202 4604 8208 4616
rect 8163 4576 8208 4604
rect 7561 4567 7619 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 9306 4604 9312 4616
rect 8435 4576 9312 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4604 10839 4607
rect 11054 4604 11060 4616
rect 10827 4576 11060 4604
rect 10827 4573 10839 4576
rect 10781 4567 10839 4573
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12618 4604 12624 4616
rect 12575 4576 12624 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12618 4564 12624 4576
rect 12676 4604 12682 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 12676 4576 13369 4604
rect 12676 4564 12682 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 13357 4567 13415 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 15105 4607 15163 4613
rect 14516 4576 14609 4604
rect 14516 4564 14522 4576
rect 15105 4573 15117 4607
rect 15151 4573 15163 4607
rect 17310 4604 17316 4616
rect 17271 4576 17316 4604
rect 15105 4567 15163 4573
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 14292 4536 14320 4564
rect 9539 4508 14320 4536
rect 14369 4539 14427 4545
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 14369 4505 14381 4539
rect 14415 4536 14427 4539
rect 15120 4536 15148 4567
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 14415 4508 15148 4536
rect 14415 4505 14427 4508
rect 14369 4499 14427 4505
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 16022 4536 16028 4548
rect 15252 4508 16028 4536
rect 15252 4496 15258 4508
rect 16022 4496 16028 4508
rect 16080 4536 16086 4548
rect 17512 4536 17540 4567
rect 17586 4564 17592 4616
rect 17644 4604 17650 4616
rect 18141 4607 18199 4613
rect 17644 4576 17689 4604
rect 17644 4564 17650 4576
rect 18141 4573 18153 4607
rect 18187 4604 18199 4607
rect 18230 4604 18236 4616
rect 18187 4576 18236 4604
rect 18187 4573 18199 4576
rect 18141 4567 18199 4573
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 16080 4508 17540 4536
rect 16080 4496 16086 4508
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 1949 4471 2007 4477
rect 1949 4468 1961 4471
rect 1728 4440 1961 4468
rect 1728 4428 1734 4440
rect 1949 4437 1961 4440
rect 1995 4437 2007 4471
rect 1949 4431 2007 4437
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5169 4471 5227 4477
rect 5169 4468 5181 4471
rect 5132 4440 5181 4468
rect 5132 4428 5138 4440
rect 5169 4437 5181 4440
rect 5215 4437 5227 4471
rect 5169 4431 5227 4437
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 9122 4468 9128 4480
rect 7892 4440 9128 4468
rect 7892 4428 7898 4440
rect 9122 4428 9128 4440
rect 9180 4468 9186 4480
rect 9401 4471 9459 4477
rect 9401 4468 9413 4471
rect 9180 4440 9413 4468
rect 9180 4428 9186 4440
rect 9401 4437 9413 4440
rect 9447 4437 9459 4471
rect 9401 4431 9459 4437
rect 13449 4471 13507 4477
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 13538 4468 13544 4480
rect 13495 4440 13544 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 15746 4468 15752 4480
rect 15519 4440 15752 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 16942 4428 16948 4480
rect 17000 4468 17006 4480
rect 17129 4471 17187 4477
rect 17129 4468 17141 4471
rect 17000 4440 17141 4468
rect 17000 4428 17006 4440
rect 17129 4437 17141 4440
rect 17175 4437 17187 4471
rect 18230 4468 18236 4480
rect 18191 4440 18236 4468
rect 17129 4431 17187 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 1104 4378 19412 4400
rect 1104 4326 7052 4378
rect 7104 4326 7116 4378
rect 7168 4326 7180 4378
rect 7232 4326 7244 4378
rect 7296 4326 7308 4378
rect 7360 4326 13155 4378
rect 13207 4326 13219 4378
rect 13271 4326 13283 4378
rect 13335 4326 13347 4378
rect 13399 4326 13411 4378
rect 13463 4326 19412 4378
rect 1104 4304 19412 4326
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 2406 4264 2412 4276
rect 2271 4236 2412 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 14277 4267 14335 4273
rect 14277 4233 14289 4267
rect 14323 4264 14335 4267
rect 14918 4264 14924 4276
rect 14323 4236 14924 4264
rect 14323 4233 14335 4236
rect 14277 4227 14335 4233
rect 14918 4224 14924 4236
rect 14976 4224 14982 4276
rect 1964 4168 2176 4196
rect 1964 4137 1992 4168
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4097 2099 4131
rect 2148 4128 2176 4168
rect 5074 4156 5080 4208
rect 5132 4156 5138 4208
rect 12710 4156 12716 4208
rect 12768 4196 12774 4208
rect 12805 4199 12863 4205
rect 12805 4196 12817 4199
rect 12768 4168 12817 4196
rect 12768 4156 12774 4168
rect 12805 4165 12817 4168
rect 12851 4165 12863 4199
rect 12805 4159 12863 4165
rect 13538 4156 13544 4208
rect 13596 4156 13602 4208
rect 16942 4196 16948 4208
rect 16903 4168 16948 4196
rect 16942 4156 16948 4168
rect 17000 4156 17006 4208
rect 18230 4196 18236 4208
rect 18170 4168 18236 4196
rect 18230 4156 18236 4168
rect 18288 4156 18294 4208
rect 3050 4128 3056 4140
rect 2148 4100 3056 4128
rect 2041 4091 2099 4097
rect 2056 4060 2084 4091
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6362 4128 6368 4140
rect 5859 4100 6368 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 8110 4128 8116 4140
rect 8071 4100 8116 4128
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 15010 4128 15016 4140
rect 14971 4100 15016 4128
rect 15010 4088 15016 4100
rect 15068 4088 15074 4140
rect 15286 4128 15292 4140
rect 15247 4100 15292 4128
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 3145 4063 3203 4069
rect 3145 4060 3157 4063
rect 2056 4032 3157 4060
rect 3145 4029 3157 4032
rect 3191 4060 3203 4063
rect 4065 4063 4123 4069
rect 4065 4060 4077 4063
rect 3191 4032 4077 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 4065 4029 4077 4032
rect 4111 4029 4123 4063
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 4065 4023 4123 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 8018 4020 8024 4072
rect 8076 4060 8082 4072
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 8076 4032 8309 4060
rect 8076 4020 8082 4032
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8297 4023 8355 4029
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14516 4032 15117 4060
rect 14516 4020 14522 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 15252 4032 15297 4060
rect 15252 4020 15258 4032
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16632 4032 16681 4060
rect 16632 4020 16638 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 2130 3952 2136 4004
rect 2188 3992 2194 4004
rect 2685 3995 2743 4001
rect 2685 3992 2697 3995
rect 2188 3964 2697 3992
rect 2188 3952 2194 3964
rect 2685 3961 2697 3964
rect 2731 3961 2743 3995
rect 2685 3955 2743 3961
rect 7374 3924 7380 3936
rect 7335 3896 7380 3924
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 7524 3896 7941 3924
rect 7524 3884 7530 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 14829 3927 14887 3933
rect 14829 3924 14841 3927
rect 14608 3896 14841 3924
rect 14608 3884 14614 3896
rect 14829 3893 14841 3896
rect 14875 3893 14887 3927
rect 14829 3887 14887 3893
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18104 3896 18429 3924
rect 18104 3884 18110 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18417 3887 18475 3893
rect 1104 3834 19412 3856
rect 1104 3782 4001 3834
rect 4053 3782 4065 3834
rect 4117 3782 4129 3834
rect 4181 3782 4193 3834
rect 4245 3782 4257 3834
rect 4309 3782 10104 3834
rect 10156 3782 10168 3834
rect 10220 3782 10232 3834
rect 10284 3782 10296 3834
rect 10348 3782 10360 3834
rect 10412 3782 16206 3834
rect 16258 3782 16270 3834
rect 16322 3782 16334 3834
rect 16386 3782 16398 3834
rect 16450 3782 16462 3834
rect 16514 3782 19412 3834
rect 1104 3760 19412 3782
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 3108 3692 3157 3720
rect 3108 3680 3114 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 3145 3683 3203 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 14921 3723 14979 3729
rect 14921 3689 14933 3723
rect 14967 3720 14979 3723
rect 15010 3720 15016 3732
rect 14967 3692 15016 3720
rect 14967 3689 14979 3692
rect 14921 3683 14979 3689
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 17681 3723 17739 3729
rect 17681 3720 17693 3723
rect 17368 3692 17693 3720
rect 17368 3680 17374 3692
rect 17681 3689 17693 3692
rect 17727 3689 17739 3723
rect 17681 3683 17739 3689
rect 7653 3655 7711 3661
rect 7653 3652 7665 3655
rect 6840 3624 7665 3652
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 1670 3584 1676 3596
rect 1631 3556 1676 3584
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 6840 3593 6868 3624
rect 7653 3621 7665 3624
rect 7699 3621 7711 3655
rect 7653 3615 7711 3621
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17770 3652 17776 3664
rect 17267 3624 17776 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17770 3612 17776 3624
rect 17828 3652 17834 3664
rect 17828 3624 18000 3652
rect 17828 3612 17834 3624
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6696 3556 6837 3584
rect 6696 3544 6702 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7101 3587 7159 3593
rect 6972 3556 7017 3584
rect 6972 3544 6978 3556
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7466 3584 7472 3596
rect 7147 3556 7472 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 8110 3584 8116 3596
rect 8023 3556 8116 3584
rect 8110 3544 8116 3556
rect 8168 3584 8174 3596
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8168 3556 8953 3584
rect 8168 3544 8174 3556
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10008 3556 10425 3584
rect 10008 3544 10014 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3584 10747 3587
rect 12526 3584 12532 3596
rect 10735 3556 12532 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 14918 3584 14924 3596
rect 14691 3556 14924 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 14918 3544 14924 3556
rect 14976 3544 14982 3596
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3584 15531 3587
rect 16482 3584 16488 3596
rect 15519 3556 16488 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 17972 3593 18000 3624
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3516 7067 3519
rect 7834 3516 7840 3528
rect 7055 3488 7840 3516
rect 7055 3485 7067 3488
rect 7009 3479 7067 3485
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 8018 3516 8024 3528
rect 7979 3488 8024 3516
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3516 14611 3519
rect 14734 3516 14740 3528
rect 14599 3488 14740 3516
rect 14599 3485 14611 3488
rect 14553 3479 14611 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 18046 3516 18052 3528
rect 18007 3488 18052 3516
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 2682 3408 2688 3460
rect 2740 3408 2746 3460
rect 9766 3408 9772 3460
rect 9824 3408 9830 3460
rect 12710 3448 12716 3460
rect 12671 3420 12716 3448
rect 12710 3408 12716 3420
rect 12768 3408 12774 3460
rect 15746 3448 15752 3460
rect 15707 3420 15752 3448
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 16206 3408 16212 3460
rect 16264 3408 16270 3460
rect 6641 3383 6699 3389
rect 6641 3349 6653 3383
rect 6687 3380 6699 3383
rect 6822 3380 6828 3392
rect 6687 3352 6828 3380
rect 6687 3349 6699 3352
rect 6641 3343 6699 3349
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 1104 3290 19412 3312
rect 1104 3238 7052 3290
rect 7104 3238 7116 3290
rect 7168 3238 7180 3290
rect 7232 3238 7244 3290
rect 7296 3238 7308 3290
rect 7360 3238 13155 3290
rect 13207 3238 13219 3290
rect 13271 3238 13283 3290
rect 13335 3238 13347 3290
rect 13399 3238 13411 3290
rect 13463 3238 19412 3290
rect 1104 3216 19412 3238
rect 2593 3179 2651 3185
rect 2593 3145 2605 3179
rect 2639 3176 2651 3179
rect 2682 3176 2688 3188
rect 2639 3148 2688 3176
rect 2639 3145 2651 3148
rect 2593 3139 2651 3145
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 8168 3148 8309 3176
rect 8168 3136 8174 3148
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 8297 3139 8355 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 14550 3176 14556 3188
rect 13280 3148 14556 3176
rect 6822 3108 6828 3120
rect 6783 3080 6828 3108
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 7374 3068 7380 3120
rect 7432 3068 7438 3120
rect 13280 3117 13308 3148
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 14734 3176 14740 3188
rect 14695 3148 14740 3176
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3176 15991 3179
rect 16206 3176 16212 3188
rect 15979 3148 16212 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 17586 3176 17592 3188
rect 17547 3148 17592 3176
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 13265 3111 13323 3117
rect 13265 3077 13277 3111
rect 13311 3077 13323 3111
rect 13265 3071 13323 3077
rect 14274 3068 14280 3120
rect 14332 3068 14338 3120
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 3418 3040 3424 3052
rect 2731 3012 3424 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 3418 3000 3424 3012
rect 3476 3000 3482 3052
rect 6362 3000 6368 3052
rect 6420 3040 6426 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6420 3012 6561 3040
rect 6420 3000 6426 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9640 3012 9873 3040
rect 9640 3000 9646 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 11112 3012 12357 3040
rect 11112 3000 11118 3012
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12584 3012 13001 3040
rect 12584 3000 12590 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 14608 3012 15853 3040
rect 14608 3000 14614 3012
rect 15841 3009 15853 3012
rect 15887 3009 15899 3043
rect 17770 3040 17776 3052
rect 17731 3012 17776 3040
rect 15841 3003 15899 3009
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 17957 3043 18015 3049
rect 17957 3009 17969 3043
rect 18003 3040 18015 3043
rect 18046 3040 18052 3052
rect 18003 3012 18052 3040
rect 18003 3009 18015 3012
rect 17957 3003 18015 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 12710 2972 12716 2984
rect 12544 2944 12716 2972
rect 12544 2913 12572 2944
rect 12710 2932 12716 2944
rect 12768 2972 12774 2984
rect 14568 2972 14596 3000
rect 12768 2944 14596 2972
rect 12768 2932 12774 2944
rect 12529 2907 12587 2913
rect 12529 2873 12541 2907
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 1104 2746 19412 2768
rect 1104 2694 4001 2746
rect 4053 2694 4065 2746
rect 4117 2694 4129 2746
rect 4181 2694 4193 2746
rect 4245 2694 4257 2746
rect 4309 2694 10104 2746
rect 10156 2694 10168 2746
rect 10220 2694 10232 2746
rect 10284 2694 10296 2746
rect 10348 2694 10360 2746
rect 10412 2694 16206 2746
rect 16258 2694 16270 2746
rect 16322 2694 16334 2746
rect 16386 2694 16398 2746
rect 16450 2694 16462 2746
rect 16514 2694 19412 2746
rect 1104 2672 19412 2694
rect 14185 2635 14243 2641
rect 14185 2601 14197 2635
rect 14231 2632 14243 2635
rect 14274 2632 14280 2644
rect 14231 2604 14280 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 10594 2564 10600 2576
rect 10555 2536 10600 2564
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2428 14335 2431
rect 14550 2428 14556 2440
rect 14323 2400 14556 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 10226 2320 10232 2372
rect 10284 2360 10290 2372
rect 10413 2363 10471 2369
rect 10413 2360 10425 2363
rect 10284 2332 10425 2360
rect 10284 2320 10290 2332
rect 10413 2329 10425 2332
rect 10459 2329 10471 2363
rect 10413 2323 10471 2329
rect 1104 2202 19412 2224
rect 1104 2150 7052 2202
rect 7104 2150 7116 2202
rect 7168 2150 7180 2202
rect 7232 2150 7244 2202
rect 7296 2150 7308 2202
rect 7360 2150 13155 2202
rect 13207 2150 13219 2202
rect 13271 2150 13283 2202
rect 13335 2150 13347 2202
rect 13399 2150 13411 2202
rect 13463 2150 19412 2202
rect 1104 2128 19412 2150
<< via1 >>
rect 4001 20102 4053 20154
rect 4065 20102 4117 20154
rect 4129 20102 4181 20154
rect 4193 20102 4245 20154
rect 4257 20102 4309 20154
rect 10104 20102 10156 20154
rect 10168 20102 10220 20154
rect 10232 20102 10284 20154
rect 10296 20102 10348 20154
rect 10360 20102 10412 20154
rect 16206 20102 16258 20154
rect 16270 20102 16322 20154
rect 16334 20102 16386 20154
rect 16398 20102 16450 20154
rect 16462 20102 16514 20154
rect 296 19864 348 19916
rect 2780 19864 2832 19916
rect 3884 19864 3936 19916
rect 6552 19907 6604 19916
rect 6552 19873 6561 19907
rect 6561 19873 6595 19907
rect 6595 19873 6604 19907
rect 6552 19864 6604 19873
rect 7104 19864 7156 19916
rect 9312 19864 9364 19916
rect 1584 19796 1636 19848
rect 3056 19839 3108 19848
rect 3056 19805 3065 19839
rect 3065 19805 3099 19839
rect 3099 19805 3108 19839
rect 3056 19796 3108 19805
rect 5448 19839 5500 19848
rect 5448 19805 5457 19839
rect 5457 19805 5491 19839
rect 5491 19805 5500 19839
rect 5448 19796 5500 19805
rect 6184 19796 6236 19848
rect 7748 19796 7800 19848
rect 8668 19796 8720 19848
rect 10416 19839 10468 19848
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 4160 19728 4212 19780
rect 7564 19728 7616 19780
rect 9864 19728 9916 19780
rect 10968 19796 11020 19848
rect 11704 19796 11756 19848
rect 20168 19932 20220 19984
rect 15752 19864 15804 19916
rect 15568 19796 15620 19848
rect 17684 19864 17736 19916
rect 18052 19907 18104 19916
rect 18052 19873 18061 19907
rect 18061 19873 18095 19907
rect 18095 19873 18104 19907
rect 18052 19864 18104 19873
rect 17132 19796 17184 19848
rect 18144 19839 18196 19848
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 11060 19728 11112 19780
rect 13636 19728 13688 19780
rect 14004 19728 14056 19780
rect 18236 19728 18288 19780
rect 4896 19660 4948 19712
rect 5080 19660 5132 19712
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 18512 19703 18564 19712
rect 18512 19669 18521 19703
rect 18521 19669 18555 19703
rect 18555 19669 18564 19703
rect 18512 19660 18564 19669
rect 7052 19558 7104 19610
rect 7116 19558 7168 19610
rect 7180 19558 7232 19610
rect 7244 19558 7296 19610
rect 7308 19558 7360 19610
rect 13155 19558 13207 19610
rect 13219 19558 13271 19610
rect 13283 19558 13335 19610
rect 13347 19558 13399 19610
rect 13411 19558 13463 19610
rect 5172 19456 5224 19508
rect 5448 19456 5500 19508
rect 10600 19456 10652 19508
rect 10968 19499 11020 19508
rect 10968 19465 10977 19499
rect 10977 19465 11011 19499
rect 11011 19465 11020 19499
rect 10968 19456 11020 19465
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 3332 19320 3384 19372
rect 4712 19320 4764 19372
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 8852 19388 8904 19440
rect 10232 19388 10284 19440
rect 6736 19320 6788 19329
rect 10692 19320 10744 19372
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 12900 19388 12952 19440
rect 16672 19456 16724 19508
rect 15200 19388 15252 19440
rect 17960 19388 18012 19440
rect 18512 19388 18564 19440
rect 10784 19320 10836 19329
rect 848 19252 900 19304
rect 2136 19252 2188 19304
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 6644 19295 6696 19304
rect 6644 19261 6653 19295
rect 6653 19261 6687 19295
rect 6687 19261 6696 19295
rect 6644 19252 6696 19261
rect 8024 19252 8076 19304
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 12440 19252 12492 19304
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 1492 19184 1544 19236
rect 4160 19184 4212 19236
rect 5816 19184 5868 19236
rect 6920 19184 6972 19236
rect 2872 19116 2924 19168
rect 3608 19116 3660 19168
rect 5540 19116 5592 19168
rect 6092 19116 6144 19168
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 15660 19159 15712 19168
rect 15660 19125 15669 19159
rect 15669 19125 15703 19159
rect 15703 19125 15712 19159
rect 15660 19116 15712 19125
rect 15844 19116 15896 19168
rect 4001 19014 4053 19066
rect 4065 19014 4117 19066
rect 4129 19014 4181 19066
rect 4193 19014 4245 19066
rect 4257 19014 4309 19066
rect 10104 19014 10156 19066
rect 10168 19014 10220 19066
rect 10232 19014 10284 19066
rect 10296 19014 10348 19066
rect 10360 19014 10412 19066
rect 16206 19014 16258 19066
rect 16270 19014 16322 19066
rect 16334 19014 16386 19066
rect 16398 19014 16450 19066
rect 16462 19014 16514 19066
rect 3056 18912 3108 18964
rect 8024 18955 8076 18964
rect 8024 18921 8033 18955
rect 8033 18921 8067 18955
rect 8067 18921 8076 18955
rect 8024 18912 8076 18921
rect 10508 18912 10560 18964
rect 14556 18912 14608 18964
rect 16028 18912 16080 18964
rect 4068 18844 4120 18896
rect 12440 18887 12492 18896
rect 12440 18853 12449 18887
rect 12449 18853 12483 18887
rect 12483 18853 12492 18887
rect 12440 18844 12492 18853
rect 5816 18819 5868 18828
rect 5816 18785 5825 18819
rect 5825 18785 5859 18819
rect 5859 18785 5868 18819
rect 5816 18776 5868 18785
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 7380 18776 7432 18828
rect 10784 18776 10836 18828
rect 12164 18819 12216 18828
rect 12164 18785 12173 18819
rect 12173 18785 12207 18819
rect 12207 18785 12216 18819
rect 12164 18776 12216 18785
rect 14556 18776 14608 18828
rect 15844 18844 15896 18896
rect 3792 18708 3844 18760
rect 3884 18708 3936 18760
rect 4068 18751 4120 18760
rect 4068 18717 4077 18751
rect 4077 18717 4111 18751
rect 4111 18717 4120 18751
rect 4068 18708 4120 18717
rect 4436 18708 4488 18760
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 8300 18708 8352 18760
rect 9404 18708 9456 18760
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 2136 18640 2188 18692
rect 2872 18683 2924 18692
rect 2872 18649 2881 18683
rect 2881 18649 2915 18683
rect 2915 18649 2924 18683
rect 2872 18640 2924 18649
rect 5724 18640 5776 18692
rect 7472 18640 7524 18692
rect 9588 18640 9640 18692
rect 12256 18708 12308 18760
rect 14280 18708 14332 18760
rect 15660 18776 15712 18828
rect 16120 18776 16172 18828
rect 17040 18776 17092 18828
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 17592 18708 17644 18760
rect 18328 18708 18380 18760
rect 3148 18572 3200 18624
rect 4344 18572 4396 18624
rect 11336 18572 11388 18624
rect 14832 18572 14884 18624
rect 7052 18470 7104 18522
rect 7116 18470 7168 18522
rect 7180 18470 7232 18522
rect 7244 18470 7296 18522
rect 7308 18470 7360 18522
rect 13155 18470 13207 18522
rect 13219 18470 13271 18522
rect 13283 18470 13335 18522
rect 13347 18470 13399 18522
rect 13411 18470 13463 18522
rect 2872 18368 2924 18420
rect 3884 18368 3936 18420
rect 4620 18368 4672 18420
rect 5080 18300 5132 18352
rect 5540 18343 5592 18352
rect 5540 18309 5549 18343
rect 5549 18309 5583 18343
rect 5583 18309 5592 18343
rect 5540 18300 5592 18309
rect 2780 18232 2832 18284
rect 3148 18275 3200 18284
rect 3148 18241 3157 18275
rect 3157 18241 3191 18275
rect 3191 18241 3200 18275
rect 3148 18232 3200 18241
rect 5816 18275 5868 18284
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 6644 18368 6696 18420
rect 8852 18368 8904 18420
rect 9956 18368 10008 18420
rect 12900 18411 12952 18420
rect 5816 18232 5868 18241
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 9128 18232 9180 18284
rect 3608 18096 3660 18148
rect 4528 18096 4580 18148
rect 6552 18164 6604 18216
rect 8208 18164 8260 18216
rect 9864 18232 9916 18284
rect 9956 18164 10008 18216
rect 6736 18096 6788 18148
rect 12900 18377 12909 18411
rect 12909 18377 12943 18411
rect 12943 18377 12952 18411
rect 12900 18368 12952 18377
rect 14188 18368 14240 18420
rect 11428 18300 11480 18352
rect 15200 18300 15252 18352
rect 18880 18368 18932 18420
rect 16580 18300 16632 18352
rect 12900 18232 12952 18284
rect 14648 18275 14700 18284
rect 14648 18241 14657 18275
rect 14657 18241 14691 18275
rect 14691 18241 14700 18275
rect 14648 18232 14700 18241
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 16672 18275 16724 18284
rect 16672 18241 16681 18275
rect 16681 18241 16715 18275
rect 16715 18241 16724 18275
rect 16672 18232 16724 18241
rect 10508 18164 10560 18216
rect 10876 18164 10928 18216
rect 11244 18164 11296 18216
rect 13912 18164 13964 18216
rect 14556 18207 14608 18216
rect 14556 18173 14565 18207
rect 14565 18173 14599 18207
rect 14599 18173 14608 18207
rect 14556 18164 14608 18173
rect 16120 18164 16172 18216
rect 16948 18207 17000 18216
rect 16948 18173 16957 18207
rect 16957 18173 16991 18207
rect 16991 18173 17000 18207
rect 16948 18164 17000 18173
rect 15200 18096 15252 18148
rect 15844 18139 15896 18148
rect 15844 18105 15853 18139
rect 15853 18105 15887 18139
rect 15887 18105 15896 18139
rect 15844 18096 15896 18105
rect 4804 18028 4856 18080
rect 10508 18028 10560 18080
rect 11152 18028 11204 18080
rect 12716 18028 12768 18080
rect 13912 18028 13964 18080
rect 15292 18028 15344 18080
rect 17040 18028 17092 18080
rect 18420 18071 18472 18080
rect 18420 18037 18429 18071
rect 18429 18037 18463 18071
rect 18463 18037 18472 18071
rect 18420 18028 18472 18037
rect 4001 17926 4053 17978
rect 4065 17926 4117 17978
rect 4129 17926 4181 17978
rect 4193 17926 4245 17978
rect 4257 17926 4309 17978
rect 10104 17926 10156 17978
rect 10168 17926 10220 17978
rect 10232 17926 10284 17978
rect 10296 17926 10348 17978
rect 10360 17926 10412 17978
rect 16206 17926 16258 17978
rect 16270 17926 16322 17978
rect 16334 17926 16386 17978
rect 16398 17926 16450 17978
rect 16462 17926 16514 17978
rect 2136 17867 2188 17876
rect 2136 17833 2145 17867
rect 2145 17833 2179 17867
rect 2179 17833 2188 17867
rect 2136 17824 2188 17833
rect 4804 17824 4856 17876
rect 16580 17824 16632 17876
rect 16948 17824 17000 17876
rect 18236 17756 18288 17808
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 5540 17688 5592 17740
rect 10692 17731 10744 17740
rect 1952 17620 2004 17672
rect 4344 17620 4396 17672
rect 4528 17663 4580 17672
rect 4528 17629 4537 17663
rect 4537 17629 4571 17663
rect 4571 17629 4580 17663
rect 4528 17620 4580 17629
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 5724 17620 5776 17672
rect 10692 17697 10701 17731
rect 10701 17697 10735 17731
rect 10735 17697 10744 17731
rect 10692 17688 10744 17697
rect 12256 17731 12308 17740
rect 12256 17697 12265 17731
rect 12265 17697 12299 17731
rect 12299 17697 12308 17731
rect 12256 17688 12308 17697
rect 15108 17688 15160 17740
rect 6920 17663 6972 17672
rect 6920 17629 6929 17663
rect 6929 17629 6963 17663
rect 6963 17629 6972 17663
rect 6920 17620 6972 17629
rect 9312 17620 9364 17672
rect 11244 17620 11296 17672
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 10508 17552 10560 17604
rect 10968 17552 11020 17604
rect 13084 17620 13136 17672
rect 13544 17620 13596 17672
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14648 17620 14700 17672
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 15936 17620 15988 17672
rect 18052 17688 18104 17740
rect 19524 17688 19576 17740
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 16120 17552 16172 17604
rect 18144 17620 18196 17672
rect 17316 17552 17368 17604
rect 3884 17484 3936 17536
rect 4436 17484 4488 17536
rect 4988 17484 5040 17536
rect 6644 17484 6696 17536
rect 7656 17484 7708 17536
rect 9680 17484 9732 17536
rect 10784 17484 10836 17536
rect 11796 17484 11848 17536
rect 14464 17484 14516 17536
rect 7052 17382 7104 17434
rect 7116 17382 7168 17434
rect 7180 17382 7232 17434
rect 7244 17382 7296 17434
rect 7308 17382 7360 17434
rect 13155 17382 13207 17434
rect 13219 17382 13271 17434
rect 13283 17382 13335 17434
rect 13347 17382 13399 17434
rect 13411 17382 13463 17434
rect 8208 17280 8260 17332
rect 9312 17280 9364 17332
rect 13544 17280 13596 17332
rect 16580 17280 16632 17332
rect 3884 17255 3936 17264
rect 3884 17221 3893 17255
rect 3893 17221 3927 17255
rect 3927 17221 3936 17255
rect 3884 17212 3936 17221
rect 6920 17212 6972 17264
rect 11796 17255 11848 17264
rect 11796 17221 11805 17255
rect 11805 17221 11839 17255
rect 11839 17221 11848 17255
rect 11796 17212 11848 17221
rect 12808 17212 12860 17264
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 4988 17144 5040 17196
rect 5816 17144 5868 17196
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 9680 17144 9732 17196
rect 10692 17144 10744 17196
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 14464 17187 14516 17196
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 15384 17144 15436 17196
rect 16948 17144 17000 17196
rect 3608 17119 3660 17128
rect 3608 17085 3617 17119
rect 3617 17085 3651 17119
rect 3651 17085 3660 17119
rect 3608 17076 3660 17085
rect 3884 17076 3936 17128
rect 6000 17076 6052 17128
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 9772 17076 9824 17085
rect 14556 17119 14608 17128
rect 14556 17085 14565 17119
rect 14565 17085 14599 17119
rect 14599 17085 14608 17119
rect 14556 17076 14608 17085
rect 18420 17144 18472 17196
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 18052 17008 18104 17060
rect 4344 16940 4396 16992
rect 10876 16940 10928 16992
rect 14740 16983 14792 16992
rect 14740 16949 14749 16983
rect 14749 16949 14783 16983
rect 14783 16949 14792 16983
rect 14740 16940 14792 16949
rect 15752 16940 15804 16992
rect 4001 16838 4053 16890
rect 4065 16838 4117 16890
rect 4129 16838 4181 16890
rect 4193 16838 4245 16890
rect 4257 16838 4309 16890
rect 10104 16838 10156 16890
rect 10168 16838 10220 16890
rect 10232 16838 10284 16890
rect 10296 16838 10348 16890
rect 10360 16838 10412 16890
rect 16206 16838 16258 16890
rect 16270 16838 16322 16890
rect 16334 16838 16386 16890
rect 16398 16838 16450 16890
rect 16462 16838 16514 16890
rect 6000 16779 6052 16788
rect 6000 16745 6009 16779
rect 6009 16745 6043 16779
rect 6043 16745 6052 16779
rect 6000 16736 6052 16745
rect 12256 16736 12308 16788
rect 5172 16668 5224 16720
rect 3608 16600 3660 16652
rect 3792 16600 3844 16652
rect 4344 16600 4396 16652
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 1860 16464 1912 16516
rect 4252 16575 4304 16584
rect 4252 16541 4261 16575
rect 4261 16541 4295 16575
rect 4295 16541 4304 16575
rect 4252 16532 4304 16541
rect 6552 16600 6604 16652
rect 5724 16575 5776 16584
rect 5724 16541 5733 16575
rect 5733 16541 5767 16575
rect 5767 16541 5776 16575
rect 5724 16532 5776 16541
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 10232 16600 10284 16652
rect 10784 16668 10836 16720
rect 12164 16668 12216 16720
rect 14740 16779 14792 16788
rect 14740 16745 14770 16779
rect 14770 16745 14792 16779
rect 14740 16736 14792 16745
rect 18236 16736 18288 16788
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 10968 16600 11020 16652
rect 12992 16643 13044 16652
rect 12992 16609 13001 16643
rect 13001 16609 13035 16643
rect 13035 16609 13044 16643
rect 12992 16600 13044 16609
rect 16672 16600 16724 16652
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 9772 16532 9824 16584
rect 12072 16532 12124 16584
rect 13544 16532 13596 16584
rect 2596 16396 2648 16448
rect 5540 16464 5592 16516
rect 6736 16464 6788 16516
rect 15752 16464 15804 16516
rect 17224 16507 17276 16516
rect 17224 16473 17233 16507
rect 17233 16473 17267 16507
rect 17267 16473 17276 16507
rect 17224 16464 17276 16473
rect 17684 16464 17736 16516
rect 8024 16396 8076 16448
rect 15384 16396 15436 16448
rect 7052 16294 7104 16346
rect 7116 16294 7168 16346
rect 7180 16294 7232 16346
rect 7244 16294 7296 16346
rect 7308 16294 7360 16346
rect 13155 16294 13207 16346
rect 13219 16294 13271 16346
rect 13283 16294 13335 16346
rect 13347 16294 13399 16346
rect 13411 16294 13463 16346
rect 1860 16235 1912 16244
rect 1860 16201 1869 16235
rect 1869 16201 1903 16235
rect 1903 16201 1912 16235
rect 1860 16192 1912 16201
rect 4252 16192 4304 16244
rect 5724 16192 5776 16244
rect 6368 16192 6420 16244
rect 1952 16099 2004 16108
rect 1952 16065 1961 16099
rect 1961 16065 1995 16099
rect 1995 16065 2004 16099
rect 1952 16056 2004 16065
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 3884 16056 3936 16108
rect 4344 16056 4396 16108
rect 4620 16056 4672 16108
rect 6644 16124 6696 16176
rect 6736 16099 6788 16108
rect 6736 16065 6746 16099
rect 6746 16065 6780 16099
rect 6780 16065 6788 16099
rect 6736 16056 6788 16065
rect 9772 16192 9824 16244
rect 12808 16192 12860 16244
rect 14648 16192 14700 16244
rect 15936 16192 15988 16244
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 17960 16192 18012 16244
rect 8024 16167 8076 16176
rect 8024 16133 8033 16167
rect 8033 16133 8067 16167
rect 8067 16133 8076 16167
rect 8024 16124 8076 16133
rect 9036 16124 9088 16176
rect 13820 16124 13872 16176
rect 10508 16056 10560 16108
rect 12900 16056 12952 16108
rect 13636 16056 13688 16108
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 15108 16124 15160 16176
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 16580 16056 16632 16108
rect 17500 16056 17552 16108
rect 2964 16031 3016 16040
rect 2964 15997 2973 16031
rect 2973 15997 3007 16031
rect 3007 15997 3016 16031
rect 2964 15988 3016 15997
rect 3976 15988 4028 16040
rect 6552 16031 6604 16040
rect 6552 15997 6561 16031
rect 6561 15997 6595 16031
rect 6595 15997 6604 16031
rect 6552 15988 6604 15997
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 6920 15988 6972 16040
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 3884 15920 3936 15972
rect 9220 15920 9272 15972
rect 16856 15920 16908 15972
rect 4344 15895 4396 15904
rect 4344 15861 4353 15895
rect 4353 15861 4387 15895
rect 4387 15861 4396 15895
rect 4344 15852 4396 15861
rect 5448 15852 5500 15904
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 4001 15750 4053 15802
rect 4065 15750 4117 15802
rect 4129 15750 4181 15802
rect 4193 15750 4245 15802
rect 4257 15750 4309 15802
rect 10104 15750 10156 15802
rect 10168 15750 10220 15802
rect 10232 15750 10284 15802
rect 10296 15750 10348 15802
rect 10360 15750 10412 15802
rect 16206 15750 16258 15802
rect 16270 15750 16322 15802
rect 16334 15750 16386 15802
rect 16398 15750 16450 15802
rect 16462 15750 16514 15802
rect 6552 15648 6604 15700
rect 9036 15691 9088 15700
rect 9036 15657 9045 15691
rect 9045 15657 9079 15691
rect 9079 15657 9088 15691
rect 9036 15648 9088 15657
rect 10508 15648 10560 15700
rect 12992 15648 13044 15700
rect 17684 15648 17736 15700
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 8116 15512 8168 15564
rect 11520 15555 11572 15564
rect 11520 15521 11529 15555
rect 11529 15521 11563 15555
rect 11563 15521 11572 15555
rect 11520 15512 11572 15521
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 4344 15444 4396 15496
rect 5172 15487 5224 15496
rect 5172 15453 5181 15487
rect 5181 15453 5215 15487
rect 5215 15453 5224 15487
rect 5172 15444 5224 15453
rect 7288 15376 7340 15428
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9956 15444 10008 15496
rect 10784 15444 10836 15496
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15844 15444 15896 15496
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 16948 15444 17000 15496
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 18236 15444 18288 15496
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 5264 15308 5316 15360
rect 7380 15308 7432 15360
rect 13360 15376 13412 15428
rect 17132 15376 17184 15428
rect 15200 15351 15252 15360
rect 15200 15317 15209 15351
rect 15209 15317 15243 15351
rect 15243 15317 15252 15351
rect 15200 15308 15252 15317
rect 16580 15308 16632 15360
rect 16764 15308 16816 15360
rect 17960 15308 18012 15360
rect 7052 15206 7104 15258
rect 7116 15206 7168 15258
rect 7180 15206 7232 15258
rect 7244 15206 7296 15258
rect 7308 15206 7360 15258
rect 13155 15206 13207 15258
rect 13219 15206 13271 15258
rect 13283 15206 13335 15258
rect 13347 15206 13399 15258
rect 13411 15206 13463 15258
rect 6920 15147 6972 15156
rect 6920 15113 6929 15147
rect 6929 15113 6963 15147
rect 6963 15113 6972 15147
rect 6920 15104 6972 15113
rect 14464 15104 14516 15156
rect 16580 15104 16632 15156
rect 16948 15104 17000 15156
rect 17316 15104 17368 15156
rect 18420 15147 18472 15156
rect 18420 15113 18429 15147
rect 18429 15113 18463 15147
rect 18463 15113 18472 15147
rect 18420 15104 18472 15113
rect 6368 15036 6420 15088
rect 1952 14968 2004 15020
rect 3884 14968 3936 15020
rect 6828 14968 6880 15020
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 7380 14968 7432 15020
rect 9036 15036 9088 15088
rect 11520 15036 11572 15088
rect 13084 15036 13136 15088
rect 9956 14968 10008 15020
rect 11152 14968 11204 15020
rect 15108 15036 15160 15088
rect 9220 14900 9272 14952
rect 14096 14968 14148 15020
rect 15200 14968 15252 15020
rect 15660 15036 15712 15088
rect 17960 15036 18012 15088
rect 15844 14968 15896 15020
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 15476 14943 15528 14952
rect 15476 14909 15485 14943
rect 15485 14909 15519 14943
rect 15519 14909 15528 14943
rect 15476 14900 15528 14909
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 14556 14832 14608 14884
rect 8116 14764 8168 14816
rect 9680 14764 9732 14816
rect 10508 14764 10560 14816
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 14004 14807 14056 14816
rect 14004 14773 14013 14807
rect 14013 14773 14047 14807
rect 14047 14773 14056 14807
rect 14004 14764 14056 14773
rect 4001 14662 4053 14714
rect 4065 14662 4117 14714
rect 4129 14662 4181 14714
rect 4193 14662 4245 14714
rect 4257 14662 4309 14714
rect 10104 14662 10156 14714
rect 10168 14662 10220 14714
rect 10232 14662 10284 14714
rect 10296 14662 10348 14714
rect 10360 14662 10412 14714
rect 16206 14662 16258 14714
rect 16270 14662 16322 14714
rect 16334 14662 16386 14714
rect 16398 14662 16450 14714
rect 16462 14662 16514 14714
rect 5080 14560 5132 14612
rect 1952 14356 2004 14408
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 2136 14288 2188 14340
rect 3608 14356 3660 14408
rect 3792 14424 3844 14476
rect 5172 14424 5224 14476
rect 6368 14560 6420 14612
rect 7472 14560 7524 14612
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 14004 14560 14056 14612
rect 15844 14603 15896 14612
rect 15844 14569 15853 14603
rect 15853 14569 15887 14603
rect 15887 14569 15896 14603
rect 15844 14560 15896 14569
rect 16948 14560 17000 14612
rect 16856 14492 16908 14544
rect 10324 14467 10376 14476
rect 3516 14288 3568 14340
rect 1952 14220 2004 14272
rect 3700 14220 3752 14272
rect 6184 14356 6236 14408
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 10324 14433 10333 14467
rect 10333 14433 10367 14467
rect 10367 14433 10376 14467
rect 10324 14424 10376 14433
rect 13452 14424 13504 14476
rect 16672 14424 16724 14476
rect 16764 14424 16816 14476
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 18236 14467 18288 14476
rect 18236 14433 18245 14467
rect 18245 14433 18279 14467
rect 18279 14433 18288 14467
rect 18236 14424 18288 14433
rect 18696 14424 18748 14476
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 10508 14356 10560 14408
rect 4528 14288 4580 14340
rect 5264 14331 5316 14340
rect 5264 14297 5273 14331
rect 5273 14297 5307 14331
rect 5307 14297 5316 14331
rect 5264 14288 5316 14297
rect 14004 14356 14056 14408
rect 16856 14399 16908 14408
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 17316 14356 17368 14408
rect 18420 14356 18472 14408
rect 4344 14220 4396 14272
rect 11428 14220 11480 14272
rect 11888 14220 11940 14272
rect 15384 14288 15436 14340
rect 13636 14220 13688 14272
rect 7052 14118 7104 14170
rect 7116 14118 7168 14170
rect 7180 14118 7232 14170
rect 7244 14118 7296 14170
rect 7308 14118 7360 14170
rect 13155 14118 13207 14170
rect 13219 14118 13271 14170
rect 13283 14118 13335 14170
rect 13347 14118 13399 14170
rect 13411 14118 13463 14170
rect 3792 14016 3844 14068
rect 3884 14016 3936 14068
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 15108 14016 15160 14068
rect 16580 14016 16632 14068
rect 17960 14016 18012 14068
rect 1952 13948 2004 14000
rect 2136 13948 2188 14000
rect 3608 13991 3660 14000
rect 3608 13957 3617 13991
rect 3617 13957 3651 13991
rect 3651 13957 3660 13991
rect 3608 13948 3660 13957
rect 8944 13948 8996 14000
rect 3700 13880 3752 13932
rect 6184 13880 6236 13932
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 9312 13880 9364 13932
rect 3148 13855 3200 13864
rect 3148 13821 3157 13855
rect 3157 13821 3191 13855
rect 3191 13821 3200 13855
rect 3148 13812 3200 13821
rect 9680 13812 9732 13864
rect 10324 13880 10376 13932
rect 11152 13948 11204 14000
rect 11428 13948 11480 14000
rect 11888 13948 11940 14000
rect 13084 13948 13136 14000
rect 10968 13880 11020 13932
rect 11060 13880 11112 13932
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 14188 13880 14240 13932
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 9864 13812 9916 13864
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 14004 13812 14056 13864
rect 14832 13812 14884 13864
rect 17040 13880 17092 13932
rect 6092 13676 6144 13728
rect 13544 13676 13596 13728
rect 4001 13574 4053 13626
rect 4065 13574 4117 13626
rect 4129 13574 4181 13626
rect 4193 13574 4245 13626
rect 4257 13574 4309 13626
rect 10104 13574 10156 13626
rect 10168 13574 10220 13626
rect 10232 13574 10284 13626
rect 10296 13574 10348 13626
rect 10360 13574 10412 13626
rect 16206 13574 16258 13626
rect 16270 13574 16322 13626
rect 16334 13574 16386 13626
rect 16398 13574 16450 13626
rect 16462 13574 16514 13626
rect 2504 13472 2556 13524
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 6828 13472 6880 13524
rect 10692 13472 10744 13524
rect 10968 13472 11020 13524
rect 3700 13336 3752 13388
rect 3148 13268 3200 13320
rect 3516 13268 3568 13320
rect 4436 13336 4488 13388
rect 4620 13268 4672 13320
rect 11336 13404 11388 13456
rect 5908 13379 5960 13388
rect 5908 13345 5917 13379
rect 5917 13345 5951 13379
rect 5951 13345 5960 13379
rect 5908 13336 5960 13345
rect 15384 13472 15436 13524
rect 18696 13515 18748 13524
rect 18696 13481 18705 13515
rect 18705 13481 18739 13515
rect 18739 13481 18748 13515
rect 18696 13472 18748 13481
rect 13452 13336 13504 13388
rect 14740 13336 14792 13388
rect 16028 13379 16080 13388
rect 7472 13268 7524 13320
rect 8392 13268 8444 13320
rect 9312 13268 9364 13320
rect 9772 13268 9824 13320
rect 10508 13268 10560 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 13636 13268 13688 13320
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 16672 13336 16724 13388
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 6920 13200 6972 13252
rect 7840 13243 7892 13252
rect 7840 13209 7849 13243
rect 7849 13209 7883 13243
rect 7883 13209 7892 13243
rect 7840 13200 7892 13209
rect 14004 13200 14056 13252
rect 2596 13132 2648 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 13912 13132 13964 13184
rect 15108 13132 15160 13184
rect 18512 13200 18564 13252
rect 7052 13030 7104 13082
rect 7116 13030 7168 13082
rect 7180 13030 7232 13082
rect 7244 13030 7296 13082
rect 7308 13030 7360 13082
rect 13155 13030 13207 13082
rect 13219 13030 13271 13082
rect 13283 13030 13335 13082
rect 13347 13030 13399 13082
rect 13411 13030 13463 13082
rect 5540 12928 5592 12980
rect 6736 12928 6788 12980
rect 7472 12971 7524 12980
rect 7472 12937 7481 12971
rect 7481 12937 7515 12971
rect 7515 12937 7524 12971
rect 7472 12928 7524 12937
rect 8944 12971 8996 12980
rect 8944 12937 8953 12971
rect 8953 12937 8987 12971
rect 8987 12937 8996 12971
rect 8944 12928 8996 12937
rect 11612 12928 11664 12980
rect 15660 12971 15712 12980
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 16120 12928 16172 12980
rect 18512 12971 18564 12980
rect 18512 12937 18521 12971
rect 18521 12937 18555 12971
rect 18555 12937 18564 12971
rect 18512 12928 18564 12937
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 3884 12792 3936 12844
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5908 12792 5960 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7656 12860 7708 12912
rect 7840 12860 7892 12912
rect 13912 12860 13964 12912
rect 14004 12860 14056 12912
rect 8208 12792 8260 12844
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 13544 12835 13596 12844
rect 2504 12767 2556 12776
rect 2504 12733 2513 12767
rect 2513 12733 2547 12767
rect 2547 12733 2556 12767
rect 2504 12724 2556 12733
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 9956 12724 10008 12776
rect 10508 12724 10560 12776
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 15108 12792 15160 12844
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 17960 12835 18012 12844
rect 17960 12801 17969 12835
rect 17969 12801 18003 12835
rect 18003 12801 18012 12835
rect 17960 12792 18012 12801
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 16764 12724 16816 12776
rect 2964 12699 3016 12708
rect 2964 12665 2973 12699
rect 2973 12665 3007 12699
rect 3007 12665 3016 12699
rect 2964 12656 3016 12665
rect 4988 12656 5040 12708
rect 4528 12588 4580 12640
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 7380 12656 7432 12708
rect 14372 12588 14424 12640
rect 4001 12486 4053 12538
rect 4065 12486 4117 12538
rect 4129 12486 4181 12538
rect 4193 12486 4245 12538
rect 4257 12486 4309 12538
rect 10104 12486 10156 12538
rect 10168 12486 10220 12538
rect 10232 12486 10284 12538
rect 10296 12486 10348 12538
rect 10360 12486 10412 12538
rect 16206 12486 16258 12538
rect 16270 12486 16322 12538
rect 16334 12486 16386 12538
rect 16398 12486 16450 12538
rect 16462 12486 16514 12538
rect 6552 12384 6604 12436
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 7380 12248 7432 12300
rect 7564 12180 7616 12232
rect 9956 12180 10008 12232
rect 11336 12384 11388 12436
rect 12716 12384 12768 12436
rect 13728 12384 13780 12436
rect 11152 12291 11204 12300
rect 11152 12257 11161 12291
rect 11161 12257 11195 12291
rect 11195 12257 11204 12291
rect 11152 12248 11204 12257
rect 14740 12248 14792 12300
rect 15660 12248 15712 12300
rect 2964 12112 3016 12164
rect 4528 12112 4580 12164
rect 6920 12112 6972 12164
rect 7840 12155 7892 12164
rect 7840 12121 7849 12155
rect 7849 12121 7883 12155
rect 7883 12121 7892 12155
rect 7840 12112 7892 12121
rect 8024 12155 8076 12164
rect 8024 12121 8033 12155
rect 8033 12121 8067 12155
rect 8067 12121 8076 12155
rect 8024 12112 8076 12121
rect 14004 12180 14056 12232
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 11060 12112 11112 12164
rect 11888 12112 11940 12164
rect 17868 12180 17920 12232
rect 17960 12112 18012 12164
rect 4712 12044 4764 12096
rect 10600 12044 10652 12096
rect 15936 12044 15988 12096
rect 7052 11942 7104 11994
rect 7116 11942 7168 11994
rect 7180 11942 7232 11994
rect 7244 11942 7296 11994
rect 7308 11942 7360 11994
rect 13155 11942 13207 11994
rect 13219 11942 13271 11994
rect 13283 11942 13335 11994
rect 13347 11942 13399 11994
rect 13411 11942 13463 11994
rect 7472 11840 7524 11892
rect 8392 11883 8444 11892
rect 8392 11849 8401 11883
rect 8401 11849 8435 11883
rect 8435 11849 8444 11883
rect 8392 11840 8444 11849
rect 4344 11772 4396 11824
rect 4988 11772 5040 11824
rect 11888 11840 11940 11892
rect 14740 11840 14792 11892
rect 9864 11815 9916 11824
rect 9864 11781 9873 11815
rect 9873 11781 9907 11815
rect 9907 11781 9916 11815
rect 9864 11772 9916 11781
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 3424 11704 3476 11756
rect 7380 11704 7432 11756
rect 12348 11704 12400 11756
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 12716 11704 12768 11756
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 7564 11636 7616 11688
rect 11060 11636 11112 11688
rect 14004 11704 14056 11756
rect 18144 11772 18196 11824
rect 14832 11704 14884 11756
rect 6460 11568 6512 11620
rect 8852 11568 8904 11620
rect 14188 11568 14240 11620
rect 16764 11704 16816 11756
rect 17960 11704 18012 11756
rect 16212 11636 16264 11688
rect 18052 11568 18104 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 16672 11500 16724 11552
rect 4001 11398 4053 11450
rect 4065 11398 4117 11450
rect 4129 11398 4181 11450
rect 4193 11398 4245 11450
rect 4257 11398 4309 11450
rect 10104 11398 10156 11450
rect 10168 11398 10220 11450
rect 10232 11398 10284 11450
rect 10296 11398 10348 11450
rect 10360 11398 10412 11450
rect 16206 11398 16258 11450
rect 16270 11398 16322 11450
rect 16334 11398 16386 11450
rect 16398 11398 16450 11450
rect 16462 11398 16514 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 7288 11296 7340 11348
rect 17868 11339 17920 11348
rect 17868 11305 17877 11339
rect 17877 11305 17911 11339
rect 17911 11305 17920 11339
rect 17868 11296 17920 11305
rect 8300 11228 8352 11280
rect 6368 11160 6420 11212
rect 6920 11160 6972 11212
rect 8024 11160 8076 11212
rect 12624 11160 12676 11212
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 16580 11160 16632 11212
rect 17960 11160 18012 11212
rect 3700 11092 3752 11144
rect 2412 11024 2464 11076
rect 2780 11024 2832 11076
rect 5724 11024 5776 11076
rect 6644 10956 6696 11008
rect 8852 11092 8904 11144
rect 9588 11092 9640 11144
rect 11704 11092 11756 11144
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12992 11092 13044 11144
rect 13544 11092 13596 11144
rect 13636 11092 13688 11144
rect 15568 11092 15620 11144
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 9956 11024 10008 11076
rect 15844 11024 15896 11076
rect 15936 11067 15988 11076
rect 15936 11033 15945 11067
rect 15945 11033 15979 11067
rect 15979 11033 15988 11067
rect 15936 11024 15988 11033
rect 16672 11024 16724 11076
rect 8024 10956 8076 11008
rect 9312 10999 9364 11008
rect 9312 10965 9321 10999
rect 9321 10965 9355 10999
rect 9355 10965 9364 10999
rect 9312 10956 9364 10965
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 15200 10956 15252 11008
rect 17316 10956 17368 11008
rect 7052 10854 7104 10906
rect 7116 10854 7168 10906
rect 7180 10854 7232 10906
rect 7244 10854 7296 10906
rect 7308 10854 7360 10906
rect 13155 10854 13207 10906
rect 13219 10854 13271 10906
rect 13283 10854 13335 10906
rect 13347 10854 13399 10906
rect 13411 10854 13463 10906
rect 6644 10752 6696 10804
rect 7380 10752 7432 10804
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 2964 10616 3016 10668
rect 3332 10616 3384 10668
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 6000 10684 6052 10736
rect 8024 10684 8076 10736
rect 8300 10727 8352 10736
rect 8300 10693 8309 10727
rect 8309 10693 8343 10727
rect 8343 10693 8352 10727
rect 8300 10684 8352 10693
rect 13544 10684 13596 10736
rect 14096 10684 14148 10736
rect 18052 10752 18104 10804
rect 9312 10659 9364 10668
rect 5448 10548 5500 10600
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 8208 10548 8260 10600
rect 8576 10591 8628 10600
rect 8576 10557 8585 10591
rect 8585 10557 8619 10591
rect 8619 10557 8628 10591
rect 8576 10548 8628 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 10692 10548 10744 10600
rect 12624 10480 12676 10532
rect 2872 10412 2924 10464
rect 4436 10412 4488 10464
rect 10876 10455 10928 10464
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 14096 10412 14148 10464
rect 15200 10616 15252 10668
rect 17960 10684 18012 10736
rect 15384 10548 15436 10600
rect 16580 10548 16632 10600
rect 16856 10548 16908 10600
rect 15476 10480 15528 10532
rect 17224 10548 17276 10600
rect 4001 10310 4053 10362
rect 4065 10310 4117 10362
rect 4129 10310 4181 10362
rect 4193 10310 4245 10362
rect 4257 10310 4309 10362
rect 10104 10310 10156 10362
rect 10168 10310 10220 10362
rect 10232 10310 10284 10362
rect 10296 10310 10348 10362
rect 10360 10310 10412 10362
rect 16206 10310 16258 10362
rect 16270 10310 16322 10362
rect 16334 10310 16386 10362
rect 16398 10310 16450 10362
rect 16462 10310 16514 10362
rect 2780 10208 2832 10260
rect 5448 10208 5500 10260
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 10876 10208 10928 10260
rect 17960 10208 18012 10260
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 3792 10140 3844 10192
rect 6920 10115 6972 10124
rect 6920 10081 6929 10115
rect 6929 10081 6963 10115
rect 6963 10081 6972 10115
rect 6920 10072 6972 10081
rect 8392 10072 8444 10124
rect 8576 10072 8628 10124
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 12900 10072 12952 10124
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3700 10004 3752 10056
rect 6000 10004 6052 10056
rect 7380 10004 7432 10056
rect 4068 9979 4120 9988
rect 4068 9945 4077 9979
rect 4077 9945 4111 9979
rect 4111 9945 4120 9979
rect 4068 9936 4120 9945
rect 4528 9936 4580 9988
rect 7840 9936 7892 9988
rect 9220 9979 9272 9988
rect 9220 9945 9229 9979
rect 9229 9945 9263 9979
rect 9263 9945 9272 9979
rect 9220 9936 9272 9945
rect 9956 9936 10008 9988
rect 12440 9936 12492 9988
rect 14004 9936 14056 9988
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 16764 10004 16816 10056
rect 16028 9936 16080 9988
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 6736 9911 6788 9920
rect 6736 9877 6745 9911
rect 6745 9877 6779 9911
rect 6779 9877 6788 9911
rect 6736 9868 6788 9877
rect 11704 9868 11756 9920
rect 14924 9868 14976 9920
rect 18144 9868 18196 9920
rect 7052 9766 7104 9818
rect 7116 9766 7168 9818
rect 7180 9766 7232 9818
rect 7244 9766 7296 9818
rect 7308 9766 7360 9818
rect 13155 9766 13207 9818
rect 13219 9766 13271 9818
rect 13283 9766 13335 9818
rect 13347 9766 13399 9818
rect 13411 9766 13463 9818
rect 1584 9664 1636 9716
rect 3700 9664 3752 9716
rect 4068 9664 4120 9716
rect 9220 9707 9272 9716
rect 9220 9673 9229 9707
rect 9229 9673 9263 9707
rect 9263 9673 9272 9707
rect 9220 9664 9272 9673
rect 15660 9707 15712 9716
rect 15660 9673 15669 9707
rect 15669 9673 15703 9707
rect 15703 9673 15712 9707
rect 15660 9664 15712 9673
rect 1492 9528 1544 9580
rect 2136 9528 2188 9580
rect 2964 9528 3016 9580
rect 3332 9528 3384 9580
rect 4436 9528 4488 9580
rect 5448 9528 5500 9580
rect 6736 9596 6788 9648
rect 7196 9596 7248 9648
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 9588 9596 9640 9648
rect 10692 9596 10744 9648
rect 14004 9596 14056 9648
rect 14740 9596 14792 9648
rect 18144 9596 18196 9648
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 2228 9324 2280 9376
rect 3792 9460 3844 9512
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 8392 9460 8444 9512
rect 9036 9460 9088 9512
rect 11704 9460 11756 9512
rect 11520 9392 11572 9444
rect 4344 9324 4396 9376
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 9404 9324 9456 9376
rect 12532 9324 12584 9376
rect 14924 9460 14976 9512
rect 15108 9460 15160 9512
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 14096 9324 14148 9376
rect 18512 9324 18564 9376
rect 4001 9222 4053 9274
rect 4065 9222 4117 9274
rect 4129 9222 4181 9274
rect 4193 9222 4245 9274
rect 4257 9222 4309 9274
rect 10104 9222 10156 9274
rect 10168 9222 10220 9274
rect 10232 9222 10284 9274
rect 10296 9222 10348 9274
rect 10360 9222 10412 9274
rect 16206 9222 16258 9274
rect 16270 9222 16322 9274
rect 16334 9222 16386 9274
rect 16398 9222 16450 9274
rect 16462 9222 16514 9274
rect 4528 9120 4580 9172
rect 6920 9120 6972 9172
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 7196 9052 7248 9104
rect 8300 8984 8352 9036
rect 5264 8916 5316 8968
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 8116 8916 8168 8968
rect 11060 8916 11112 8968
rect 14832 9120 14884 9172
rect 15384 9120 15436 9172
rect 17132 9120 17184 9172
rect 15844 9052 15896 9104
rect 16580 8984 16632 9036
rect 17592 8984 17644 9036
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 15108 8959 15160 8968
rect 15108 8925 15117 8959
rect 15117 8925 15151 8959
rect 15151 8925 15160 8959
rect 15108 8916 15160 8925
rect 15568 8916 15620 8968
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 3700 8848 3752 8900
rect 6092 8848 6144 8900
rect 13820 8848 13872 8900
rect 16028 8848 16080 8900
rect 18696 8916 18748 8968
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 11060 8780 11112 8832
rect 12348 8780 12400 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 14372 8780 14424 8832
rect 7052 8678 7104 8730
rect 7116 8678 7168 8730
rect 7180 8678 7232 8730
rect 7244 8678 7296 8730
rect 7308 8678 7360 8730
rect 13155 8678 13207 8730
rect 13219 8678 13271 8730
rect 13283 8678 13335 8730
rect 13347 8678 13399 8730
rect 13411 8678 13463 8730
rect 6460 8576 6512 8628
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 7564 8576 7616 8628
rect 3240 8508 3292 8560
rect 5540 8508 5592 8560
rect 1676 8440 1728 8492
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 2688 8440 2740 8492
rect 1492 8372 1544 8424
rect 3148 8483 3200 8492
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 6184 8440 6236 8492
rect 3240 8372 3292 8424
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 5448 8347 5500 8356
rect 5448 8313 5457 8347
rect 5457 8313 5491 8347
rect 5491 8313 5500 8347
rect 5448 8304 5500 8313
rect 8116 8440 8168 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 12808 8508 12860 8560
rect 14372 8576 14424 8628
rect 15384 8576 15436 8628
rect 14280 8508 14332 8560
rect 8208 8440 8260 8449
rect 8668 8440 8720 8492
rect 11060 8440 11112 8492
rect 15200 8440 15252 8492
rect 16580 8440 16632 8492
rect 18512 8440 18564 8492
rect 8300 8372 8352 8424
rect 12716 8372 12768 8424
rect 17132 8415 17184 8424
rect 9956 8304 10008 8356
rect 11244 8304 11296 8356
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 18696 8372 18748 8424
rect 1676 8236 1728 8288
rect 8760 8236 8812 8288
rect 12900 8236 12952 8288
rect 13728 8304 13780 8356
rect 14096 8304 14148 8356
rect 16948 8236 17000 8288
rect 4001 8134 4053 8186
rect 4065 8134 4117 8186
rect 4129 8134 4181 8186
rect 4193 8134 4245 8186
rect 4257 8134 4309 8186
rect 10104 8134 10156 8186
rect 10168 8134 10220 8186
rect 10232 8134 10284 8186
rect 10296 8134 10348 8186
rect 10360 8134 10412 8186
rect 16206 8134 16258 8186
rect 16270 8134 16322 8186
rect 16334 8134 16386 8186
rect 16398 8134 16450 8186
rect 16462 8134 16514 8186
rect 6368 8032 6420 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 6460 7964 6512 8016
rect 8300 8032 8352 8084
rect 12808 8032 12860 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 8944 7939 8996 7948
rect 3332 7760 3384 7812
rect 6092 7828 6144 7880
rect 7380 7828 7432 7880
rect 6184 7760 6236 7812
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 5264 7692 5316 7744
rect 6000 7735 6052 7744
rect 6000 7701 6009 7735
rect 6009 7701 6043 7735
rect 6043 7701 6052 7735
rect 6000 7692 6052 7701
rect 6644 7692 6696 7744
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 12624 7939 12676 7948
rect 12624 7905 12633 7939
rect 12633 7905 12667 7939
rect 12667 7905 12676 7939
rect 12624 7896 12676 7905
rect 12900 7939 12952 7948
rect 12900 7905 12909 7939
rect 12909 7905 12943 7939
rect 12943 7905 12952 7939
rect 12900 7896 12952 7905
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 15384 7896 15436 7948
rect 7748 7871 7800 7880
rect 7748 7837 7758 7871
rect 7758 7837 7792 7871
rect 7792 7837 7800 7871
rect 7748 7828 7800 7837
rect 12992 7828 13044 7880
rect 15476 7828 15528 7880
rect 18144 7828 18196 7880
rect 9128 7760 9180 7812
rect 10600 7760 10652 7812
rect 11244 7760 11296 7812
rect 9036 7692 9088 7744
rect 10876 7692 10928 7744
rect 18236 7692 18288 7744
rect 7052 7590 7104 7642
rect 7116 7590 7168 7642
rect 7180 7590 7232 7642
rect 7244 7590 7296 7642
rect 7308 7590 7360 7642
rect 13155 7590 13207 7642
rect 13219 7590 13271 7642
rect 13283 7590 13335 7642
rect 13347 7590 13399 7642
rect 13411 7590 13463 7642
rect 3332 7531 3384 7540
rect 3332 7497 3341 7531
rect 3341 7497 3375 7531
rect 3375 7497 3384 7531
rect 3332 7488 3384 7497
rect 6000 7488 6052 7540
rect 9128 7531 9180 7540
rect 6644 7463 6696 7472
rect 6644 7429 6653 7463
rect 6653 7429 6687 7463
rect 6687 7429 6696 7463
rect 6644 7420 6696 7429
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 10600 7488 10652 7540
rect 14740 7488 14792 7540
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 9588 7420 9640 7472
rect 3148 7352 3200 7404
rect 8760 7395 8812 7404
rect 2044 7284 2096 7336
rect 3240 7284 3292 7336
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 7380 7284 7432 7336
rect 12716 7352 12768 7404
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13820 7395 13872 7404
rect 13084 7352 13136 7361
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 10968 7284 11020 7336
rect 15016 7352 15068 7404
rect 18144 7488 18196 7540
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 18236 7420 18288 7472
rect 16764 7284 16816 7336
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 3424 7148 3476 7200
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 12992 7216 13044 7268
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 15016 7148 15068 7200
rect 4001 7046 4053 7098
rect 4065 7046 4117 7098
rect 4129 7046 4181 7098
rect 4193 7046 4245 7098
rect 4257 7046 4309 7098
rect 10104 7046 10156 7098
rect 10168 7046 10220 7098
rect 10232 7046 10284 7098
rect 10296 7046 10348 7098
rect 10360 7046 10412 7098
rect 16206 7046 16258 7098
rect 16270 7046 16322 7098
rect 16334 7046 16386 7098
rect 16398 7046 16450 7098
rect 16462 7046 16514 7098
rect 7380 6987 7432 6996
rect 7380 6953 7389 6987
rect 7389 6953 7423 6987
rect 7423 6953 7432 6987
rect 7380 6944 7432 6953
rect 9588 6987 9640 6996
rect 9588 6953 9597 6987
rect 9597 6953 9631 6987
rect 9631 6953 9640 6987
rect 9588 6944 9640 6953
rect 1400 6808 1452 6860
rect 3700 6808 3752 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 12716 6851 12768 6860
rect 12440 6808 12492 6817
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 16120 6876 16172 6928
rect 17224 6919 17276 6928
rect 16028 6851 16080 6860
rect 16028 6817 16037 6851
rect 16037 6817 16071 6851
rect 16071 6817 16080 6851
rect 17224 6885 17233 6919
rect 17233 6885 17267 6919
rect 17267 6885 17276 6919
rect 17224 6876 17276 6885
rect 16028 6808 16080 6817
rect 8116 6740 8168 6792
rect 9956 6740 10008 6792
rect 13084 6740 13136 6792
rect 15016 6740 15068 6792
rect 4068 6715 4120 6724
rect 4068 6681 4077 6715
rect 4077 6681 4111 6715
rect 4111 6681 4120 6715
rect 4068 6672 4120 6681
rect 6460 6672 6512 6724
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 16672 6740 16724 6792
rect 17316 6740 17368 6792
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 18328 6740 18380 6792
rect 7052 6502 7104 6554
rect 7116 6502 7168 6554
rect 7180 6502 7232 6554
rect 7244 6502 7296 6554
rect 7308 6502 7360 6554
rect 13155 6502 13207 6554
rect 13219 6502 13271 6554
rect 13283 6502 13335 6554
rect 13347 6502 13399 6554
rect 13411 6502 13463 6554
rect 4068 6400 4120 6452
rect 4160 6400 4212 6452
rect 4344 6400 4396 6452
rect 4896 6400 4948 6452
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 7748 6400 7800 6452
rect 13084 6400 13136 6452
rect 2688 6332 2740 6384
rect 15660 6400 15712 6452
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 2136 6264 2188 6316
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 14924 6332 14976 6384
rect 15752 6332 15804 6384
rect 5540 6264 5592 6316
rect 7840 6307 7892 6316
rect 5080 6196 5132 6248
rect 5448 6196 5500 6248
rect 4436 6128 4488 6180
rect 5264 6128 5316 6180
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 8116 6264 8168 6316
rect 12900 6264 12952 6316
rect 13728 6264 13780 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 17684 6307 17736 6316
rect 17684 6273 17693 6307
rect 17693 6273 17727 6307
rect 17727 6273 17736 6307
rect 17684 6264 17736 6273
rect 1860 6060 1912 6112
rect 12348 6196 12400 6248
rect 15568 6196 15620 6248
rect 12532 6060 12584 6112
rect 17408 6060 17460 6112
rect 4001 5958 4053 6010
rect 4065 5958 4117 6010
rect 4129 5958 4181 6010
rect 4193 5958 4245 6010
rect 4257 5958 4309 6010
rect 10104 5958 10156 6010
rect 10168 5958 10220 6010
rect 10232 5958 10284 6010
rect 10296 5958 10348 6010
rect 10360 5958 10412 6010
rect 16206 5958 16258 6010
rect 16270 5958 16322 6010
rect 16334 5958 16386 6010
rect 16398 5958 16450 6010
rect 16462 5958 16514 6010
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 7840 5856 7892 5908
rect 12348 5899 12400 5908
rect 12348 5865 12357 5899
rect 12357 5865 12391 5899
rect 12391 5865 12400 5899
rect 12348 5856 12400 5865
rect 16120 5856 16172 5908
rect 16856 5856 16908 5908
rect 2136 5720 2188 5772
rect 1400 5652 1452 5704
rect 5540 5720 5592 5772
rect 12716 5788 12768 5840
rect 9312 5720 9364 5772
rect 12440 5720 12492 5772
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 4344 5652 4396 5704
rect 5356 5652 5408 5704
rect 6368 5652 6420 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 10876 5695 10928 5704
rect 1768 5627 1820 5636
rect 1768 5593 1777 5627
rect 1777 5593 1811 5627
rect 1811 5593 1820 5627
rect 1768 5584 1820 5593
rect 3516 5584 3568 5636
rect 6920 5584 6972 5636
rect 7564 5584 7616 5636
rect 9128 5584 9180 5636
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 15568 5695 15620 5704
rect 12716 5652 12768 5661
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 16580 5652 16632 5704
rect 16948 5695 17000 5704
rect 16948 5661 16957 5695
rect 16957 5661 16991 5695
rect 16991 5661 17000 5695
rect 16948 5652 17000 5661
rect 18328 5652 18380 5704
rect 17224 5627 17276 5636
rect 17224 5593 17233 5627
rect 17233 5593 17267 5627
rect 17267 5593 17276 5627
rect 17224 5584 17276 5593
rect 4252 5516 4304 5568
rect 9404 5516 9456 5568
rect 13544 5516 13596 5568
rect 15936 5516 15988 5568
rect 7052 5414 7104 5466
rect 7116 5414 7168 5466
rect 7180 5414 7232 5466
rect 7244 5414 7296 5466
rect 7308 5414 7360 5466
rect 13155 5414 13207 5466
rect 13219 5414 13271 5466
rect 13283 5414 13335 5466
rect 13347 5414 13399 5466
rect 13411 5414 13463 5466
rect 1768 5312 1820 5364
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 11060 5312 11112 5364
rect 17224 5312 17276 5364
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 5264 5244 5316 5296
rect 9404 5287 9456 5296
rect 9404 5253 9413 5287
rect 9413 5253 9447 5287
rect 9447 5253 9456 5287
rect 9404 5244 9456 5253
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 2136 5108 2188 5160
rect 4436 5108 4488 5160
rect 7012 5176 7064 5228
rect 7656 5176 7708 5228
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 8944 5176 8996 5228
rect 8208 5108 8260 5160
rect 9496 5108 9548 5160
rect 9772 5108 9824 5160
rect 12440 5108 12492 5160
rect 13544 5176 13596 5228
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 18236 5219 18288 5228
rect 18236 5185 18245 5219
rect 18245 5185 18279 5219
rect 18279 5185 18288 5219
rect 18236 5176 18288 5185
rect 14280 5108 14332 5160
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 5540 5040 5592 5092
rect 12716 5083 12768 5092
rect 12716 5049 12725 5083
rect 12725 5049 12759 5083
rect 12759 5049 12768 5083
rect 12716 5040 12768 5049
rect 6552 4972 6604 5024
rect 9956 4972 10008 5024
rect 15292 4972 15344 5024
rect 4001 4870 4053 4922
rect 4065 4870 4117 4922
rect 4129 4870 4181 4922
rect 4193 4870 4245 4922
rect 4257 4870 4309 4922
rect 10104 4870 10156 4922
rect 10168 4870 10220 4922
rect 10232 4870 10284 4922
rect 10296 4870 10348 4922
rect 10360 4870 10412 4922
rect 16206 4870 16258 4922
rect 16270 4870 16322 4922
rect 16334 4870 16386 4922
rect 16398 4870 16450 4922
rect 16462 4870 16514 4922
rect 7564 4768 7616 4820
rect 8300 4811 8352 4820
rect 8300 4777 8309 4811
rect 8309 4777 8343 4811
rect 8343 4777 8352 4811
rect 8300 4768 8352 4777
rect 9496 4768 9548 4820
rect 12900 4768 12952 4820
rect 6920 4743 6972 4752
rect 6920 4709 6929 4743
rect 6929 4709 6963 4743
rect 6963 4709 6972 4743
rect 6920 4700 6972 4709
rect 17500 4700 17552 4752
rect 1676 4632 1728 4684
rect 2688 4632 2740 4684
rect 6644 4675 6696 4684
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 5264 4607 5316 4616
rect 2412 4564 2464 4573
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7472 4564 7524 4616
rect 9588 4632 9640 4684
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 13912 4632 13964 4684
rect 15016 4675 15068 4684
rect 15016 4641 15025 4675
rect 15025 4641 15059 4675
rect 15059 4641 15068 4675
rect 15016 4632 15068 4641
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 9312 4564 9364 4616
rect 11060 4564 11112 4616
rect 12624 4564 12676 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 15200 4496 15252 4548
rect 16028 4496 16080 4548
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 18236 4564 18288 4616
rect 1676 4428 1728 4480
rect 5080 4428 5132 4480
rect 7840 4428 7892 4480
rect 9128 4428 9180 4480
rect 13544 4428 13596 4480
rect 15752 4428 15804 4480
rect 16948 4428 17000 4480
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 7052 4326 7104 4378
rect 7116 4326 7168 4378
rect 7180 4326 7232 4378
rect 7244 4326 7296 4378
rect 7308 4326 7360 4378
rect 13155 4326 13207 4378
rect 13219 4326 13271 4378
rect 13283 4326 13335 4378
rect 13347 4326 13399 4378
rect 13411 4326 13463 4378
rect 2412 4224 2464 4276
rect 14924 4224 14976 4276
rect 5080 4156 5132 4208
rect 12716 4156 12768 4208
rect 13544 4156 13596 4208
rect 16948 4199 17000 4208
rect 16948 4165 16957 4199
rect 16957 4165 16991 4199
rect 16991 4165 17000 4199
rect 16948 4156 17000 4165
rect 18236 4156 18288 4208
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 6368 4088 6420 4140
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 15016 4131 15068 4140
rect 15016 4097 15025 4131
rect 15025 4097 15059 4131
rect 15059 4097 15068 4131
rect 15016 4088 15068 4097
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 8024 4020 8076 4072
rect 14464 4020 14516 4072
rect 15200 4063 15252 4072
rect 15200 4029 15209 4063
rect 15209 4029 15243 4063
rect 15243 4029 15252 4063
rect 15200 4020 15252 4029
rect 16580 4020 16632 4072
rect 2136 3952 2188 4004
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 7472 3884 7524 3936
rect 14556 3884 14608 3936
rect 18052 3884 18104 3936
rect 4001 3782 4053 3834
rect 4065 3782 4117 3834
rect 4129 3782 4181 3834
rect 4193 3782 4245 3834
rect 4257 3782 4309 3834
rect 10104 3782 10156 3834
rect 10168 3782 10220 3834
rect 10232 3782 10284 3834
rect 10296 3782 10348 3834
rect 10360 3782 10412 3834
rect 16206 3782 16258 3834
rect 16270 3782 16322 3834
rect 16334 3782 16386 3834
rect 16398 3782 16450 3834
rect 16462 3782 16514 3834
rect 3056 3680 3108 3732
rect 12992 3723 13044 3732
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 15016 3680 15068 3732
rect 17316 3680 17368 3732
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 6644 3544 6696 3596
rect 17776 3612 17828 3664
rect 6920 3587 6972 3596
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 7472 3544 7524 3596
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 9956 3544 10008 3596
rect 12532 3544 12584 3596
rect 14924 3544 14976 3596
rect 16488 3544 16540 3596
rect 7840 3476 7892 3528
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 14740 3476 14792 3528
rect 18052 3519 18104 3528
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 2688 3408 2740 3460
rect 9772 3408 9824 3460
rect 12716 3451 12768 3460
rect 12716 3417 12725 3451
rect 12725 3417 12759 3451
rect 12759 3417 12768 3451
rect 12716 3408 12768 3417
rect 15752 3451 15804 3460
rect 15752 3417 15761 3451
rect 15761 3417 15795 3451
rect 15795 3417 15804 3451
rect 15752 3408 15804 3417
rect 16212 3408 16264 3460
rect 6828 3340 6880 3392
rect 7052 3238 7104 3290
rect 7116 3238 7168 3290
rect 7180 3238 7232 3290
rect 7244 3238 7296 3290
rect 7308 3238 7360 3290
rect 13155 3238 13207 3290
rect 13219 3238 13271 3290
rect 13283 3238 13335 3290
rect 13347 3238 13399 3290
rect 13411 3238 13463 3290
rect 2688 3136 2740 3188
rect 8116 3136 8168 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 6828 3111 6880 3120
rect 6828 3077 6837 3111
rect 6837 3077 6871 3111
rect 6871 3077 6880 3111
rect 6828 3068 6880 3077
rect 7380 3068 7432 3120
rect 14556 3136 14608 3188
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 16212 3136 16264 3188
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 14280 3068 14332 3120
rect 3424 3000 3476 3052
rect 6368 3000 6420 3052
rect 9588 3000 9640 3052
rect 11060 3000 11112 3052
rect 12532 3000 12584 3052
rect 14556 3000 14608 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 18052 3000 18104 3052
rect 12716 2932 12768 2984
rect 4001 2694 4053 2746
rect 4065 2694 4117 2746
rect 4129 2694 4181 2746
rect 4193 2694 4245 2746
rect 4257 2694 4309 2746
rect 10104 2694 10156 2746
rect 10168 2694 10220 2746
rect 10232 2694 10284 2746
rect 10296 2694 10348 2746
rect 10360 2694 10412 2746
rect 16206 2694 16258 2746
rect 16270 2694 16322 2746
rect 16334 2694 16386 2746
rect 16398 2694 16450 2746
rect 16462 2694 16514 2746
rect 14280 2592 14332 2644
rect 10600 2567 10652 2576
rect 10600 2533 10609 2567
rect 10609 2533 10643 2567
rect 10643 2533 10652 2567
rect 10600 2524 10652 2533
rect 14556 2388 14608 2440
rect 10232 2320 10284 2372
rect 7052 2150 7104 2202
rect 7116 2150 7168 2202
rect 7180 2150 7232 2202
rect 7244 2150 7296 2202
rect 7308 2150 7360 2202
rect 13155 2150 13207 2202
rect 13219 2150 13271 2202
rect 13283 2150 13335 2202
rect 13347 2150 13399 2202
rect 13411 2150 13463 2202
<< metal2 >>
rect 294 21861 350 22661
rect 846 21861 902 22661
rect 1490 21861 1546 22661
rect 2134 21861 2190 22661
rect 2778 21861 2834 22661
rect 3330 21978 3386 22661
rect 2976 21950 3386 21978
rect 308 19922 336 21861
rect 296 19916 348 19922
rect 296 19858 348 19864
rect 860 19310 888 21861
rect 848 19304 900 19310
rect 848 19246 900 19252
rect 1504 19242 1532 21861
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1492 19236 1544 19242
rect 1492 19178 1544 19184
rect 1596 16574 1624 19790
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1504 16546 1624 16574
rect 1688 16574 1716 19314
rect 2148 19310 2176 21861
rect 2792 20074 2820 21861
rect 2792 20046 2912 20074
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2136 18692 2188 18698
rect 2136 18634 2188 18640
rect 2148 17882 2176 18634
rect 2792 18290 2820 19858
rect 2884 19174 2912 20046
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2872 18692 2924 18698
rect 2872 18634 2924 18640
rect 2884 18426 2912 18634
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 2792 17746 2820 18226
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1688 16546 1808 16574
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11354 1440 11698
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1504 9586 1532 16546
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11393 1624 11494
rect 1582 11384 1638 11393
rect 1582 11319 1638 11328
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9722 1624 9998
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1504 8430 1532 9522
rect 1688 8498 1716 10066
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1676 8288 1728 8294
rect 1676 8230 1728 8236
rect 1688 7954 1716 8230
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 6866 1440 7822
rect 1780 6914 1808 16546
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 1872 16250 1900 16458
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1964 16114 1992 17614
rect 2976 17202 3004 21950
rect 3330 21861 3386 21950
rect 3974 21861 4030 22661
rect 4618 21861 4674 22661
rect 5262 21861 5318 22661
rect 5814 21861 5870 22661
rect 6458 21978 6514 22661
rect 6458 21950 6592 21978
rect 6458 21861 6514 21950
rect 3988 20346 4016 21861
rect 3804 20318 4016 20346
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3068 18970 3096 19790
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3160 18290 3188 18566
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2608 16114 2636 16390
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 1964 15026 1992 16050
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2976 15570 3004 15982
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1964 14414 1992 14962
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1964 14006 1992 14214
rect 2148 14006 2176 14282
rect 1952 14000 2004 14006
rect 1952 13942 2004 13948
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2516 13530 2544 14350
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2516 12782 2544 13466
rect 3160 13326 3188 13806
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12850 2636 13126
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2976 12170 3004 12650
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11082 2452 11494
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10266 2820 11018
rect 3344 10674 3372 19314
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18154 3648 19110
rect 3804 18766 3832 20318
rect 4001 20156 4309 20176
rect 4001 20154 4007 20156
rect 4063 20154 4087 20156
rect 4143 20154 4167 20156
rect 4223 20154 4247 20156
rect 4303 20154 4309 20156
rect 4063 20102 4065 20154
rect 4245 20102 4247 20154
rect 4001 20100 4007 20102
rect 4063 20100 4087 20102
rect 4143 20100 4167 20102
rect 4223 20100 4247 20102
rect 4303 20100 4309 20102
rect 4001 20080 4309 20100
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3896 18766 3924 19858
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 4172 19242 4200 19722
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4001 19068 4309 19088
rect 4001 19066 4007 19068
rect 4063 19066 4087 19068
rect 4143 19066 4167 19068
rect 4223 19066 4247 19068
rect 4303 19066 4309 19068
rect 4063 19014 4065 19066
rect 4245 19014 4247 19066
rect 4001 19012 4007 19014
rect 4063 19012 4087 19014
rect 4143 19012 4167 19014
rect 4223 19012 4247 19014
rect 4303 19012 4309 19014
rect 4001 18992 4309 19012
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 4080 18766 4108 18838
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 3896 18426 3924 18702
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 4001 17980 4309 18000
rect 4001 17978 4007 17980
rect 4063 17978 4087 17980
rect 4143 17978 4167 17980
rect 4223 17978 4247 17980
rect 4303 17978 4309 17980
rect 4063 17926 4065 17978
rect 4245 17926 4247 17978
rect 4001 17924 4007 17926
rect 4063 17924 4087 17926
rect 4143 17924 4167 17926
rect 4223 17924 4247 17926
rect 4303 17924 4309 17926
rect 4001 17904 4309 17924
rect 4356 17678 4384 18566
rect 4448 18306 4476 18702
rect 4632 18426 4660 21861
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4724 18306 4752 19314
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4448 18278 4752 18306
rect 4528 18148 4580 18154
rect 4528 18090 4580 18096
rect 4540 17678 4568 18090
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 3896 17270 3924 17478
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3620 16658 3648 17070
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3804 14482 3832 16594
rect 3896 16114 3924 17070
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4001 16892 4309 16912
rect 4001 16890 4007 16892
rect 4063 16890 4087 16892
rect 4143 16890 4167 16892
rect 4223 16890 4247 16892
rect 4303 16890 4309 16892
rect 4063 16838 4065 16890
rect 4245 16838 4247 16890
rect 4001 16836 4007 16838
rect 4063 16836 4087 16838
rect 4143 16836 4167 16838
rect 4223 16836 4247 16838
rect 4303 16836 4309 16838
rect 4001 16816 4309 16836
rect 4356 16658 4384 16934
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3896 15978 3924 16050
rect 3988 16046 4016 16526
rect 4264 16250 4292 16526
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4356 16114 4384 16594
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4001 15804 4309 15824
rect 4001 15802 4007 15804
rect 4063 15802 4087 15804
rect 4143 15802 4167 15804
rect 4223 15802 4247 15804
rect 4303 15802 4309 15804
rect 4063 15750 4065 15802
rect 4245 15750 4247 15802
rect 4001 15748 4007 15750
rect 4063 15748 4087 15750
rect 4143 15748 4167 15750
rect 4223 15748 4247 15750
rect 4303 15748 4309 15750
rect 4001 15728 4309 15748
rect 4356 15502 4384 15846
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3528 13326 3556 14282
rect 3620 14006 3648 14350
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3712 13938 3740 14214
rect 3804 14074 3832 14418
rect 3896 14074 3924 14962
rect 4001 14716 4309 14736
rect 4001 14714 4007 14716
rect 4063 14714 4087 14716
rect 4143 14714 4167 14716
rect 4223 14714 4247 14716
rect 4303 14714 4309 14716
rect 4063 14662 4065 14714
rect 4245 14662 4247 14714
rect 4001 14660 4007 14662
rect 4063 14660 4087 14662
rect 4143 14660 4167 14662
rect 4223 14660 4247 14662
rect 4303 14660 4309 14662
rect 4001 14640 4309 14660
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3712 13394 3740 13874
rect 3700 13388 3752 13394
rect 3700 13330 3752 13336
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3804 12306 3832 14010
rect 3896 12850 3924 14010
rect 4001 13628 4309 13648
rect 4001 13626 4007 13628
rect 4063 13626 4087 13628
rect 4143 13626 4167 13628
rect 4223 13626 4247 13628
rect 4303 13626 4309 13628
rect 4063 13574 4065 13626
rect 4245 13574 4247 13626
rect 4001 13572 4007 13574
rect 4063 13572 4087 13574
rect 4143 13572 4167 13574
rect 4223 13572 4247 13574
rect 4303 13572 4309 13574
rect 4001 13552 4309 13572
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 4001 12540 4309 12560
rect 4001 12538 4007 12540
rect 4063 12538 4087 12540
rect 4143 12538 4167 12540
rect 4223 12538 4247 12540
rect 4303 12538 4309 12540
rect 4063 12486 4065 12538
rect 4245 12486 4247 12538
rect 4001 12484 4007 12486
rect 4063 12484 4087 12486
rect 4143 12484 4167 12486
rect 4223 12484 4247 12486
rect 4303 12484 4309 12486
rect 4001 12464 4309 12484
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 4356 11830 4384 14214
rect 4448 13394 4476 17478
rect 4632 16114 4660 18278
rect 4816 18086 4844 18702
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4816 17882 4844 18022
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14346 4568 14758
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4632 13326 4660 16050
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4540 12170 4568 12582
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2884 10062 2912 10406
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2976 9586 3004 10610
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 7342 2084 8434
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 1688 6886 1808 6914
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 5710 1440 6802
rect 1688 6322 1716 6886
rect 2148 6322 2176 9522
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 8498 2268 9318
rect 3252 8566 3280 9862
rect 3344 9586 3372 10610
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 2700 6390 2728 8434
rect 3160 7750 3188 8434
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 7410 3188 7686
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3252 7342 3280 8366
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3344 7546 3372 7754
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 3602 1440 5646
rect 1688 4690 1716 6258
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1780 5370 1808 5578
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1872 5234 1900 6054
rect 2148 5778 2176 6258
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 2148 4622 2176 5102
rect 2700 4690 2728 6326
rect 3252 5914 3280 7278
rect 3436 7206 3464 11698
rect 4001 11452 4309 11472
rect 4001 11450 4007 11452
rect 4063 11450 4087 11452
rect 4143 11450 4167 11452
rect 4223 11450 4247 11452
rect 4303 11450 4309 11452
rect 4063 11398 4065 11450
rect 4245 11398 4247 11450
rect 4001 11396 4007 11398
rect 4063 11396 4087 11398
rect 4143 11396 4167 11398
rect 4223 11396 4247 11398
rect 4303 11396 4309 11398
rect 4001 11376 4309 11396
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3712 10062 3740 11086
rect 4001 10364 4309 10384
rect 4001 10362 4007 10364
rect 4063 10362 4087 10364
rect 4143 10362 4167 10364
rect 4223 10362 4247 10364
rect 4303 10362 4309 10364
rect 4063 10310 4065 10362
rect 4245 10310 4247 10362
rect 4001 10308 4007 10310
rect 4063 10308 4087 10310
rect 4143 10308 4167 10310
rect 4223 10308 4247 10310
rect 4303 10308 4309 10310
rect 4001 10288 4309 10308
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3712 9722 3740 9998
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3712 8906 3740 9658
rect 3804 9518 3832 10134
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 4080 9722 4108 9930
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 4356 9382 4384 11766
rect 4724 10674 4752 12038
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4724 10554 4752 10610
rect 4724 10526 4844 10554
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 9586 4476 10406
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4001 9276 4309 9296
rect 4001 9274 4007 9276
rect 4063 9274 4087 9276
rect 4143 9274 4167 9276
rect 4223 9274 4247 9276
rect 4303 9274 4309 9276
rect 4063 9222 4065 9274
rect 4245 9222 4247 9274
rect 4001 9220 4007 9222
rect 4063 9220 4087 9222
rect 4143 9220 4167 9222
rect 4223 9220 4247 9222
rect 4303 9220 4309 9222
rect 4001 9200 4309 9220
rect 4540 9178 4568 9930
rect 4816 9518 4844 10526
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3712 8430 3740 8842
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 3602 1716 4422
rect 2148 4010 2176 4558
rect 2424 4282 2452 4558
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 3068 3738 3096 4082
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2700 3194 2728 3402
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 3436 3058 3464 7142
rect 3712 6866 3740 8366
rect 4001 8188 4309 8208
rect 4001 8186 4007 8188
rect 4063 8186 4087 8188
rect 4143 8186 4167 8188
rect 4223 8186 4247 8188
rect 4303 8186 4309 8188
rect 4063 8134 4065 8186
rect 4245 8134 4247 8186
rect 4001 8132 4007 8134
rect 4063 8132 4087 8134
rect 4143 8132 4167 8134
rect 4223 8132 4247 8134
rect 4303 8132 4309 8134
rect 4001 8112 4309 8132
rect 4001 7100 4309 7120
rect 4001 7098 4007 7100
rect 4063 7098 4087 7100
rect 4143 7098 4167 7100
rect 4223 7098 4247 7100
rect 4303 7098 4309 7100
rect 4063 7046 4065 7098
rect 4245 7046 4247 7098
rect 4001 7044 4007 7046
rect 4063 7044 4087 7046
rect 4143 7044 4167 7046
rect 4223 7044 4247 7046
rect 4303 7044 4309 7046
rect 4001 7024 4309 7044
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 4080 6458 4108 6666
rect 4908 6458 4936 19654
rect 5092 18358 5120 19654
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5080 18352 5132 18358
rect 5080 18294 5132 18300
rect 5184 17678 5212 19450
rect 5276 18068 5304 21861
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5460 19514 5488 19790
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5828 19242 5856 21861
rect 6564 19922 6592 21950
rect 7102 21861 7158 22661
rect 7746 21861 7802 22661
rect 8298 21861 8354 22661
rect 8942 21978 8998 22661
rect 8942 21950 9352 21978
rect 8942 21861 8998 21950
rect 7116 19922 7144 21861
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7760 19854 7788 21861
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 5552 18358 5580 19110
rect 6104 18834 6132 19110
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5276 18040 5580 18068
rect 5552 17746 5580 18040
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5736 17678 5764 18634
rect 5828 18290 5856 18770
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17202 5028 17478
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 5184 16726 5212 17614
rect 5828 17202 5856 18226
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 6012 16794 6040 17070
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 5184 15586 5212 16662
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5092 15558 5212 15586
rect 5460 15570 5488 15846
rect 5448 15564 5500 15570
rect 5092 14618 5120 15558
rect 5448 15506 5500 15512
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5184 14822 5212 15438
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5184 14482 5212 14758
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5276 14346 5304 15302
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5552 12986 5580 16458
rect 5736 16250 5764 16526
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 6196 16130 6224 19790
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7052 19612 7360 19632
rect 7052 19610 7058 19612
rect 7114 19610 7138 19612
rect 7194 19610 7218 19612
rect 7274 19610 7298 19612
rect 7354 19610 7360 19612
rect 7114 19558 7116 19610
rect 7296 19558 7298 19610
rect 7052 19556 7058 19558
rect 7114 19556 7138 19558
rect 7194 19556 7218 19558
rect 7274 19556 7298 19558
rect 7354 19556 7360 19558
rect 7052 19536 7360 19556
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6564 18222 6592 19246
rect 6656 18426 6684 19246
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6748 18154 6776 19314
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6380 16250 6408 17138
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6012 16102 6224 16130
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5920 12850 5948 13330
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5000 12714 5028 12786
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 5000 11830 5028 12650
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11082 5764 11494
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 6012 10742 6040 16102
rect 6380 15094 6408 16186
rect 6564 16046 6592 16594
rect 6656 16182 6684 17478
rect 6748 16522 6776 18090
rect 6932 17678 6960 19178
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7052 18524 7360 18544
rect 7052 18522 7058 18524
rect 7114 18522 7138 18524
rect 7194 18522 7218 18524
rect 7274 18522 7298 18524
rect 7354 18522 7360 18524
rect 7114 18470 7116 18522
rect 7296 18470 7298 18522
rect 7052 18468 7058 18470
rect 7114 18468 7138 18470
rect 7194 18468 7218 18470
rect 7274 18468 7298 18470
rect 7354 18468 7360 18470
rect 7052 18448 7360 18468
rect 7392 18290 7420 18770
rect 7484 18698 7512 19110
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 7052 17436 7360 17456
rect 7052 17434 7058 17436
rect 7114 17434 7138 17436
rect 7194 17434 7218 17436
rect 7274 17434 7298 17436
rect 7354 17434 7360 17436
rect 7114 17382 7116 17434
rect 7296 17382 7298 17434
rect 7052 17380 7058 17382
rect 7114 17380 7138 17382
rect 7194 17380 7218 17382
rect 7274 17380 7298 17382
rect 7354 17380 7360 17382
rect 7052 17360 7360 17380
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 6932 16590 6960 17206
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6656 16046 6684 16118
rect 6748 16114 6776 16458
rect 7052 16348 7360 16368
rect 7052 16346 7058 16348
rect 7114 16346 7138 16348
rect 7194 16346 7218 16348
rect 7274 16346 7298 16348
rect 7354 16346 7360 16348
rect 7114 16294 7116 16346
rect 7296 16294 7298 16346
rect 7052 16292 7058 16294
rect 7114 16292 7138 16294
rect 7194 16292 7218 16294
rect 7274 16292 7298 16294
rect 7354 16292 7360 16294
rect 7052 16272 7360 16292
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6564 15706 6592 15982
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6932 15162 6960 15982
rect 7300 15434 7512 15450
rect 7288 15428 7512 15434
rect 7340 15422 7512 15428
rect 7288 15370 7340 15376
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7052 15260 7360 15280
rect 7052 15258 7058 15260
rect 7114 15258 7138 15260
rect 7194 15258 7218 15260
rect 7274 15258 7298 15260
rect 7354 15258 7360 15260
rect 7114 15206 7116 15258
rect 7296 15206 7298 15258
rect 7052 15204 7058 15206
rect 7114 15204 7138 15206
rect 7194 15204 7218 15206
rect 7274 15204 7298 15206
rect 7354 15204 7360 15206
rect 7052 15184 7360 15204
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 6380 14618 6408 15030
rect 7392 15026 7420 15302
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13938 6224 14350
rect 6380 13938 6408 14554
rect 6840 14414 6868 14962
rect 7484 14618 7512 15422
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 13530 6132 13670
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5460 10266 5488 10542
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5460 9586 5488 10202
rect 6012 10062 6040 10678
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 7750 5304 8910
rect 6104 8906 6132 9862
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 8566 5580 8774
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4172 6322 4200 6394
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4001 6012 4309 6032
rect 4001 6010 4007 6012
rect 4063 6010 4087 6012
rect 4143 6010 4167 6012
rect 4223 6010 4247 6012
rect 4303 6010 4309 6012
rect 4063 5958 4065 6010
rect 4245 5958 4247 6010
rect 4001 5956 4007 5958
rect 4063 5956 4087 5958
rect 4143 5956 4167 5958
rect 4223 5956 4247 5958
rect 4303 5956 4309 5958
rect 4001 5936 4309 5956
rect 4356 5710 4384 6394
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3528 5370 3556 5578
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 4264 5234 4292 5510
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4448 5166 4476 6122
rect 5092 5914 5120 6190
rect 5276 6186 5304 7686
rect 5460 6254 5488 8298
rect 6104 7886 6132 8842
rect 6196 8498 6224 13874
rect 6840 13530 6868 14350
rect 7052 14172 7360 14192
rect 7052 14170 7058 14172
rect 7114 14170 7138 14172
rect 7194 14170 7218 14172
rect 7274 14170 7298 14172
rect 7354 14170 7360 14172
rect 7114 14118 7116 14170
rect 7296 14118 7298 14170
rect 7052 14116 7058 14118
rect 7114 14116 7138 14118
rect 7194 14116 7218 14118
rect 7274 14116 7298 14118
rect 7354 14116 7360 14118
rect 7052 14096 7360 14116
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 11218 6408 12582
rect 6564 12442 6592 12786
rect 6748 12782 6776 12922
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6932 12170 6960 13194
rect 7052 13084 7360 13104
rect 7052 13082 7058 13084
rect 7114 13082 7138 13084
rect 7194 13082 7218 13084
rect 7274 13082 7298 13084
rect 7354 13082 7360 13084
rect 7114 13030 7116 13082
rect 7296 13030 7298 13082
rect 7052 13028 7058 13030
rect 7114 13028 7138 13030
rect 7194 13028 7218 13030
rect 7274 13028 7298 13030
rect 7354 13028 7360 13030
rect 7052 13008 7360 13028
rect 7484 12986 7512 13262
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7392 12434 7420 12650
rect 7576 12434 7604 19722
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 8036 18970 8064 19246
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8312 18766 8340 21861
rect 9324 19922 9352 21950
rect 9586 21861 9642 22661
rect 10230 21861 10286 22661
rect 10782 21861 10838 22661
rect 11426 21861 11482 22661
rect 12070 21861 12126 22661
rect 12714 21861 12770 22661
rect 13266 21978 13322 22661
rect 13266 21950 13768 21978
rect 13266 21861 13322 21950
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8220 18222 8248 18702
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 12918 7696 17478
rect 8220 17338 8248 18158
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 8036 16182 8064 16390
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 14822 8156 15506
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14074 8156 14758
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7852 12918 7880 13194
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7392 12406 7512 12434
rect 7576 12406 7696 12434
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 7052 11996 7360 12016
rect 7052 11994 7058 11996
rect 7114 11994 7138 11996
rect 7194 11994 7218 11996
rect 7274 11994 7298 11996
rect 7354 11994 7360 11996
rect 7114 11942 7116 11994
rect 7296 11942 7298 11994
rect 7052 11940 7058 11942
rect 7114 11940 7138 11942
rect 7194 11940 7218 11942
rect 7274 11940 7298 11942
rect 7354 11940 7360 11942
rect 7052 11920 7360 11940
rect 7392 11762 7420 12242
rect 7484 11898 7512 12406
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6472 8974 6500 11562
rect 7300 11354 7328 11630
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10810 6684 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6932 10130 6960 11154
rect 7052 10908 7360 10928
rect 7052 10906 7058 10908
rect 7114 10906 7138 10908
rect 7194 10906 7218 10908
rect 7274 10906 7298 10908
rect 7354 10906 7360 10908
rect 7114 10854 7116 10906
rect 7296 10854 7298 10906
rect 7052 10852 7058 10854
rect 7114 10852 7138 10854
rect 7194 10852 7218 10854
rect 7274 10852 7298 10854
rect 7354 10852 7360 10854
rect 7052 10832 7360 10852
rect 7392 10810 7420 11698
rect 7576 11694 7604 12174
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9654 6776 9862
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6932 9178 6960 10066
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7052 9820 7360 9840
rect 7052 9818 7058 9820
rect 7114 9818 7138 9820
rect 7194 9818 7218 9820
rect 7274 9818 7298 9820
rect 7354 9818 7360 9820
rect 7114 9766 7116 9818
rect 7296 9766 7298 9818
rect 7052 9764 7058 9766
rect 7114 9764 7138 9766
rect 7194 9764 7218 9766
rect 7274 9764 7298 9766
rect 7354 9764 7360 9766
rect 7052 9744 7360 9764
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7208 9110 7236 9590
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 8634 6500 8910
rect 7052 8732 7360 8752
rect 7052 8730 7058 8732
rect 7114 8730 7138 8732
rect 7194 8730 7218 8732
rect 7274 8730 7298 8732
rect 7354 8730 7360 8732
rect 7114 8678 7116 8730
rect 7296 8678 7298 8730
rect 7052 8676 7058 8678
rect 7114 8676 7138 8678
rect 7194 8676 7218 8678
rect 7274 8676 7298 8678
rect 7354 8676 7360 8678
rect 7052 8656 7360 8676
rect 7392 8634 7420 9998
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6196 7818 6224 8434
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7546 6040 7686
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6380 7342 6408 8026
rect 6472 8022 6500 8570
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 7576 7954 7604 8570
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7478 6684 7686
rect 7052 7644 7360 7664
rect 7052 7642 7058 7644
rect 7114 7642 7138 7644
rect 7194 7642 7218 7644
rect 7274 7642 7298 7644
rect 7354 7642 7360 7644
rect 7114 7590 7116 7642
rect 7296 7590 7298 7642
rect 7052 7588 7058 7590
rect 7114 7588 7138 7590
rect 7194 7588 7218 7590
rect 7274 7588 7298 7590
rect 7354 7588 7360 7590
rect 7052 7568 7360 7588
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 7392 7342 7420 7822
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6322 5580 6598
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5276 5302 5304 6122
rect 5356 5704 5408 5710
rect 5460 5692 5488 6190
rect 5552 5778 5580 6258
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 6380 5710 6408 7278
rect 7392 7002 7420 7278
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6472 6458 6500 6666
rect 7052 6556 7360 6576
rect 7052 6554 7058 6556
rect 7114 6554 7138 6556
rect 7194 6554 7218 6556
rect 7274 6554 7298 6556
rect 7354 6554 7360 6556
rect 7114 6502 7116 6554
rect 7296 6502 7298 6554
rect 7052 6500 7058 6502
rect 7114 6500 7138 6502
rect 7194 6500 7218 6502
rect 7274 6500 7298 6502
rect 7354 6500 7360 6502
rect 7052 6480 7360 6500
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 5408 5664 5488 5692
rect 6368 5704 6420 5710
rect 5356 5646 5408 5652
rect 6368 5646 6420 5652
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4001 4924 4309 4944
rect 4001 4922 4007 4924
rect 4063 4922 4087 4924
rect 4143 4922 4167 4924
rect 4223 4922 4247 4924
rect 4303 4922 4309 4924
rect 4063 4870 4065 4922
rect 4245 4870 4247 4922
rect 4001 4868 4007 4870
rect 4063 4868 4087 4870
rect 4143 4868 4167 4870
rect 4223 4868 4247 4870
rect 4303 4868 4309 4870
rect 4001 4848 4309 4868
rect 5276 4622 5304 5238
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5092 4214 5120 4422
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5552 4078 5580 5034
rect 6380 4146 6408 5646
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4622 6592 4966
rect 6932 4758 6960 5578
rect 7052 5468 7360 5488
rect 7052 5466 7058 5468
rect 7114 5466 7138 5468
rect 7194 5466 7218 5468
rect 7274 5466 7298 5468
rect 7354 5466 7360 5468
rect 7114 5414 7116 5466
rect 7296 5414 7298 5466
rect 7052 5412 7058 5414
rect 7114 5412 7138 5414
rect 7194 5412 7218 5414
rect 7274 5412 7298 5414
rect 7354 5412 7360 5414
rect 7052 5392 7360 5412
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 4001 3836 4309 3856
rect 4001 3834 4007 3836
rect 4063 3834 4087 3836
rect 4143 3834 4167 3836
rect 4223 3834 4247 3836
rect 4303 3834 4309 3836
rect 4063 3782 4065 3834
rect 4245 3782 4247 3834
rect 4001 3780 4007 3782
rect 4063 3780 4087 3782
rect 4143 3780 4167 3782
rect 4223 3780 4247 3782
rect 4303 3780 4309 3782
rect 4001 3760 4309 3780
rect 6380 3058 6408 4082
rect 6656 3602 6684 4626
rect 7024 4604 7052 5170
rect 7576 4826 7604 5578
rect 7668 5234 7696 12406
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7852 9994 7880 12106
rect 8036 11218 8064 12106
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8036 10742 8064 10950
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 8220 10606 8248 12786
rect 8404 11898 8432 13262
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8312 10742 8340 11222
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 8974 8156 9318
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8128 8498 8156 8910
rect 8220 8498 8248 10542
rect 8588 10130 8616 10542
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8404 9518 8432 10066
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 6458 7788 7822
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7852 6322 7880 6802
rect 8128 6798 8156 7142
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 6322 8156 6734
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7852 5914 7880 6258
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 8220 5166 8248 8434
rect 8312 8430 8340 8978
rect 8680 8498 8708 19790
rect 8852 19440 8904 19446
rect 8852 19382 8904 19388
rect 8864 18426 8892 19382
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9140 17202 9168 18226
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9324 17338 9352 17614
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9048 15706 9076 16118
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9140 15502 9168 17138
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 9048 14618 9076 15030
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9140 14414 9168 15438
rect 9232 14958 9260 15914
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 12986 8984 13942
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9324 13326 9352 13874
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 11626 8892 12786
rect 9416 12434 9444 18702
rect 9600 18698 9628 21861
rect 10244 20346 10272 21861
rect 9968 20318 10272 20346
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9876 18290 9904 19722
rect 9968 18426 9996 20318
rect 10104 20156 10412 20176
rect 10104 20154 10110 20156
rect 10166 20154 10190 20156
rect 10246 20154 10270 20156
rect 10326 20154 10350 20156
rect 10406 20154 10412 20156
rect 10166 20102 10168 20154
rect 10348 20102 10350 20154
rect 10104 20100 10110 20102
rect 10166 20100 10190 20102
rect 10246 20100 10270 20102
rect 10326 20100 10350 20102
rect 10406 20100 10412 20102
rect 10104 20080 10412 20100
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10244 19446 10272 19654
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10428 19258 10456 19790
rect 10796 19530 10824 21861
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10600 19508 10652 19514
rect 10796 19502 10916 19530
rect 10980 19514 11008 19790
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 10600 19450 10652 19456
rect 10612 19310 10640 19450
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10600 19304 10652 19310
rect 10428 19230 10548 19258
rect 10600 19246 10652 19252
rect 10104 19068 10412 19088
rect 10104 19066 10110 19068
rect 10166 19066 10190 19068
rect 10246 19066 10270 19068
rect 10326 19066 10350 19068
rect 10406 19066 10412 19068
rect 10166 19014 10168 19066
rect 10348 19014 10350 19066
rect 10104 19012 10110 19014
rect 10166 19012 10190 19014
rect 10246 19012 10270 19014
rect 10326 19012 10350 19014
rect 10406 19012 10412 19014
rect 10104 18992 10412 19012
rect 10520 18970 10548 19230
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 10520 18222 10548 18906
rect 10612 18766 10640 19246
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17202 9720 17478
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 16658 9720 17138
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9784 16590 9812 17070
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9784 16250 9812 16526
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9968 15502 9996 18158
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10104 17980 10412 18000
rect 10104 17978 10110 17980
rect 10166 17978 10190 17980
rect 10246 17978 10270 17980
rect 10326 17978 10350 17980
rect 10406 17978 10412 17980
rect 10166 17926 10168 17978
rect 10348 17926 10350 17978
rect 10104 17924 10110 17926
rect 10166 17924 10190 17926
rect 10246 17924 10270 17926
rect 10326 17924 10350 17926
rect 10406 17924 10412 17926
rect 10104 17904 10412 17924
rect 10520 17610 10548 18022
rect 10704 17746 10732 19314
rect 10796 18834 10824 19314
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10888 18222 10916 19502
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11072 19394 11100 19722
rect 10980 19366 11100 19394
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10704 17202 10732 17682
rect 10980 17610 11008 19366
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10104 16892 10412 16912
rect 10104 16890 10110 16892
rect 10166 16890 10190 16892
rect 10246 16890 10270 16892
rect 10326 16890 10350 16892
rect 10406 16890 10412 16892
rect 10166 16838 10168 16890
rect 10348 16838 10350 16890
rect 10104 16836 10110 16838
rect 10166 16836 10190 16838
rect 10246 16836 10270 16838
rect 10326 16836 10350 16838
rect 10406 16836 10412 16838
rect 10104 16816 10412 16836
rect 10796 16726 10824 17478
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10244 16046 10272 16594
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10104 15804 10412 15824
rect 10104 15802 10110 15804
rect 10166 15802 10190 15804
rect 10246 15802 10270 15804
rect 10326 15802 10350 15804
rect 10406 15802 10412 15804
rect 10166 15750 10168 15802
rect 10348 15750 10350 15802
rect 10104 15748 10110 15750
rect 10166 15748 10190 15750
rect 10246 15748 10270 15750
rect 10326 15748 10350 15750
rect 10406 15748 10412 15750
rect 10104 15728 10412 15748
rect 10520 15706 10548 16050
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10796 15502 10824 16662
rect 10888 16658 10916 16934
rect 10980 16658 11008 17546
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 9968 15026 9996 15438
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 13870 9720 14758
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9692 13410 9720 13806
rect 9692 13382 9812 13410
rect 9784 13326 9812 13382
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9416 12406 9536 12434
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11150 8892 11562
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10674 9352 10950
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 8090 8340 8366
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8772 7410 8800 8230
rect 8956 7954 8984 10066
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 9722 9260 9930
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9416 9586 9444 10542
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8956 5234 8984 7890
rect 9048 7750 9076 9454
rect 9416 9382 9444 9522
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 5624 9076 7686
rect 9140 7546 9168 7754
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9508 5794 9536 12406
rect 9876 11830 9904 13806
rect 9968 12782 9996 14962
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10104 14716 10412 14736
rect 10104 14714 10110 14716
rect 10166 14714 10190 14716
rect 10246 14714 10270 14716
rect 10326 14714 10350 14716
rect 10406 14714 10412 14716
rect 10166 14662 10168 14714
rect 10348 14662 10350 14714
rect 10104 14660 10110 14662
rect 10166 14660 10190 14662
rect 10246 14660 10270 14662
rect 10326 14660 10350 14662
rect 10406 14660 10412 14662
rect 10104 14640 10412 14660
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 13938 10364 14418
rect 10520 14414 10548 14758
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10980 13938 11008 16594
rect 11164 15026 11192 18022
rect 11256 17678 11284 18158
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11164 14006 11192 14962
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10104 13628 10412 13648
rect 10104 13626 10110 13628
rect 10166 13626 10190 13628
rect 10246 13626 10270 13628
rect 10326 13626 10350 13628
rect 10406 13626 10412 13628
rect 10166 13574 10168 13626
rect 10348 13574 10350 13626
rect 10104 13572 10110 13574
rect 10166 13572 10190 13574
rect 10246 13572 10270 13574
rect 10326 13572 10350 13574
rect 10406 13572 10412 13574
rect 10104 13552 10412 13572
rect 10704 13530 10732 13806
rect 10980 13530 11008 13874
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10520 12782 10548 13262
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 9968 12238 9996 12718
rect 10104 12540 10412 12560
rect 10104 12538 10110 12540
rect 10166 12538 10190 12540
rect 10246 12538 10270 12540
rect 10326 12538 10350 12540
rect 10406 12538 10412 12540
rect 10166 12486 10168 12538
rect 10348 12486 10350 12538
rect 10104 12484 10110 12486
rect 10166 12484 10190 12486
rect 10246 12484 10270 12486
rect 10326 12484 10350 12486
rect 10406 12484 10412 12486
rect 10104 12464 10412 12484
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9600 9654 9628 11086
rect 9968 11082 9996 12174
rect 10104 11452 10412 11472
rect 10104 11450 10110 11452
rect 10166 11450 10190 11452
rect 10246 11450 10270 11452
rect 10326 11450 10350 11452
rect 10406 11450 10412 11452
rect 10166 11398 10168 11450
rect 10348 11398 10350 11450
rect 10104 11396 10110 11398
rect 10166 11396 10190 11398
rect 10246 11396 10270 11398
rect 10326 11396 10350 11398
rect 10406 11396 10412 11398
rect 10104 11376 10412 11396
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 10520 10606 10548 12718
rect 11072 12170 11100 13874
rect 11348 13462 11376 18566
rect 11440 18358 11468 21861
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11532 15570 11560 17138
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11532 15094 11560 15506
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11440 14006 11468 14214
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11532 13938 11560 15030
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12306 11192 13126
rect 11348 12442 11376 13398
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12986 11652 13262
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 10674 10640 12038
rect 11072 11694 11100 12106
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11716 11150 11744 19790
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11808 17270 11836 17478
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 12084 16590 12112 21861
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12452 18902 12480 19246
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12176 17678 12204 18770
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12268 17746 12296 18702
rect 12728 18086 12756 21861
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13155 19612 13463 19632
rect 13155 19610 13161 19612
rect 13217 19610 13241 19612
rect 13297 19610 13321 19612
rect 13377 19610 13401 19612
rect 13457 19610 13463 19612
rect 13217 19558 13219 19610
rect 13399 19558 13401 19610
rect 13155 19556 13161 19558
rect 13217 19556 13241 19558
rect 13297 19556 13321 19558
rect 13377 19556 13401 19558
rect 13457 19556 13463 19558
rect 13155 19536 13463 19556
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 12912 18426 12940 19382
rect 13155 18524 13463 18544
rect 13155 18522 13161 18524
rect 13217 18522 13241 18524
rect 13297 18522 13321 18524
rect 13377 18522 13401 18524
rect 13457 18522 13463 18524
rect 13217 18470 13219 18522
rect 13399 18470 13401 18522
rect 13155 18468 13161 18470
rect 13217 18468 13241 18470
rect 13297 18468 13321 18470
rect 13377 18468 13401 18470
rect 13457 18468 13463 18470
rect 13155 18448 13463 18468
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 16726 12204 17614
rect 12268 16794 12296 17682
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12820 16250 12848 17206
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12912 16114 12940 18226
rect 13084 17672 13136 17678
rect 13004 17632 13084 17660
rect 13004 16658 13032 17632
rect 13084 17614 13136 17620
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13155 17436 13463 17456
rect 13155 17434 13161 17436
rect 13217 17434 13241 17436
rect 13297 17434 13321 17436
rect 13377 17434 13401 17436
rect 13457 17434 13463 17436
rect 13217 17382 13219 17434
rect 13399 17382 13401 17434
rect 13155 17380 13161 17382
rect 13217 17380 13241 17382
rect 13297 17380 13321 17382
rect 13377 17380 13401 17382
rect 13457 17380 13463 17382
rect 13155 17360 13463 17380
rect 13556 17338 13584 17614
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 13004 15706 13032 16594
rect 13556 16590 13584 17274
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13155 16348 13463 16368
rect 13155 16346 13161 16348
rect 13217 16346 13241 16348
rect 13297 16346 13321 16348
rect 13377 16346 13401 16348
rect 13457 16346 13463 16348
rect 13217 16294 13219 16346
rect 13399 16294 13401 16346
rect 13155 16292 13161 16294
rect 13217 16292 13241 16294
rect 13297 16292 13321 16294
rect 13377 16292 13401 16294
rect 13457 16292 13463 16294
rect 13155 16272 13463 16292
rect 13648 16266 13676 19722
rect 13740 18034 13768 21950
rect 13910 21861 13966 22661
rect 14554 21861 14610 22661
rect 15198 21861 15254 22661
rect 15750 21861 15806 22661
rect 16394 21978 16450 22661
rect 16132 21950 16450 21978
rect 13924 18222 13952 21861
rect 14004 19780 14056 19786
rect 14004 19722 14056 19728
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13912 18080 13964 18086
rect 13740 18006 13860 18034
rect 13912 18022 13964 18028
rect 13556 16238 13676 16266
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13372 15434 13400 15846
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13155 15260 13463 15280
rect 13155 15258 13161 15260
rect 13217 15258 13241 15260
rect 13297 15258 13321 15260
rect 13377 15258 13401 15260
rect 13457 15258 13463 15260
rect 13217 15206 13219 15258
rect 13399 15206 13401 15258
rect 13155 15204 13161 15206
rect 13217 15204 13241 15206
rect 13297 15204 13321 15206
rect 13377 15204 13401 15206
rect 13457 15204 13463 15206
rect 13155 15184 13463 15204
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 14006 11928 14214
rect 13096 14006 13124 15030
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14482 13492 14758
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13155 14172 13463 14192
rect 13155 14170 13161 14172
rect 13217 14170 13241 14172
rect 13297 14170 13321 14172
rect 13377 14170 13401 14172
rect 13457 14170 13463 14172
rect 13217 14118 13219 14170
rect 13399 14118 13401 14170
rect 13155 14116 13161 14118
rect 13217 14116 13241 14118
rect 13297 14116 13321 14118
rect 13377 14116 13401 14118
rect 13457 14116 13463 14118
rect 13155 14096 13463 14116
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13556 13818 13584 16238
rect 13832 16182 13860 18006
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13924 16114 13952 18022
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13648 14278 13676 16050
rect 14016 15994 14044 19722
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14200 18426 14228 19246
rect 14568 18970 14596 21861
rect 15212 19530 15240 21861
rect 15764 19922 15792 21861
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15212 19502 15332 19530
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14292 17678 14320 18702
rect 14568 18222 14596 18770
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 18290 14872 18566
rect 15212 18358 15240 19382
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14476 17202 14504 17478
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14568 17134 14596 18158
rect 14660 17678 14688 18226
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14660 16250 14688 17614
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 16794 14780 16934
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 15120 16182 15148 17682
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 13832 15966 14044 15994
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13464 13790 13584 13818
rect 13464 13394 13492 13790
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13155 13084 13463 13104
rect 13155 13082 13161 13084
rect 13217 13082 13241 13084
rect 13297 13082 13321 13084
rect 13377 13082 13401 13084
rect 13457 13082 13463 13084
rect 13217 13030 13219 13082
rect 13399 13030 13401 13082
rect 13155 13028 13161 13030
rect 13217 13028 13241 13030
rect 13297 13028 13321 13030
rect 13377 13028 13401 13030
rect 13457 13028 13463 13030
rect 13155 13008 13463 13028
rect 13556 12850 13584 13670
rect 13648 13326 13676 14214
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 12728 12442 12756 12786
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13740 12442 13768 12718
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 13728 12436 13780 12442
rect 13832 12434 13860 15966
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14108 15026 14136 15846
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14476 15162 14504 15438
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14568 14890 14596 15506
rect 15120 15094 15148 16118
rect 15212 16114 15240 18090
rect 15304 18086 15332 19502
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15396 17202 15424 17614
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15396 15502 15424 16390
rect 15384 15496 15436 15502
rect 15436 15444 15516 15450
rect 15384 15438 15516 15444
rect 15396 15422 15516 15438
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 14618 14044 14758
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14016 13870 14044 14350
rect 15120 14074 15148 15030
rect 15212 15026 15240 15302
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15488 14958 15516 15422
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12918 13952 13126
rect 14016 12918 14044 13194
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 13832 12406 13952 12434
rect 13728 12378 13780 12384
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11900 11898 11928 12106
rect 13155 11996 13463 12016
rect 13155 11994 13161 11996
rect 13217 11994 13241 11996
rect 13297 11994 13321 11996
rect 13377 11994 13401 11996
rect 13457 11994 13463 11996
rect 13217 11942 13219 11994
rect 13399 11942 13401 11994
rect 13155 11940 13161 11942
rect 13217 11940 13241 11942
rect 13297 11940 13321 11942
rect 13377 11940 13401 11942
rect 13457 11940 13463 11942
rect 13155 11920 13463 11940
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12360 11150 12388 11698
rect 12636 11218 12664 11698
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10104 10364 10412 10384
rect 10104 10362 10110 10364
rect 10166 10362 10190 10364
rect 10246 10362 10270 10364
rect 10326 10362 10350 10364
rect 10406 10362 10412 10364
rect 10166 10310 10168 10362
rect 10348 10310 10350 10362
rect 10104 10308 10110 10310
rect 10166 10308 10190 10310
rect 10246 10308 10270 10310
rect 10326 10308 10350 10310
rect 10406 10308 10412 10310
rect 10104 10288 10412 10308
rect 10704 10266 10732 10542
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 10888 10266 10916 10406
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9968 9178 9996 9930
rect 10704 9654 10732 10202
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 11532 9450 11560 10406
rect 11716 9926 11744 10610
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9518 11744 9862
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 10104 9276 10412 9296
rect 10104 9274 10110 9276
rect 10166 9274 10190 9276
rect 10246 9274 10270 9276
rect 10326 9274 10350 9276
rect 10406 9274 10412 9276
rect 10166 9222 10168 9274
rect 10348 9222 10350 9274
rect 10104 9220 10110 9222
rect 10166 9220 10190 9222
rect 10246 9220 10270 9222
rect 10326 9220 10350 9222
rect 10406 9220 10412 9222
rect 10104 9200 10412 9220
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8838 11100 8910
rect 12360 8838 12388 11086
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 9994 12480 10950
rect 12728 10810 12756 11698
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11150 13676 11494
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 11072 8498 11100 8774
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 9968 7546 9996 8298
rect 10104 8188 10412 8208
rect 10104 8186 10110 8188
rect 10166 8186 10190 8188
rect 10246 8186 10270 8188
rect 10326 8186 10350 8188
rect 10406 8186 10412 8188
rect 10166 8134 10168 8186
rect 10348 8134 10350 8186
rect 10104 8132 10110 8134
rect 10166 8132 10190 8134
rect 10246 8132 10270 8134
rect 10326 8132 10350 8134
rect 10406 8132 10412 8134
rect 10104 8112 10412 8132
rect 11256 7818 11284 8298
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 10612 7546 10640 7754
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9600 7002 9628 7414
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9324 5778 9536 5794
rect 9312 5772 9536 5778
rect 9364 5766 9536 5772
rect 9312 5714 9364 5720
rect 9128 5636 9180 5642
rect 9048 5596 9128 5624
rect 9128 5578 9180 5584
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 8220 4622 8248 5102
rect 8312 4826 8340 5170
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 6932 4576 7052 4604
rect 7472 4616 7524 4622
rect 6932 3602 6960 4576
rect 7472 4558 7524 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7052 4380 7360 4400
rect 7052 4378 7058 4380
rect 7114 4378 7138 4380
rect 7194 4378 7218 4380
rect 7274 4378 7298 4380
rect 7354 4378 7360 4380
rect 7114 4326 7116 4378
rect 7296 4326 7298 4378
rect 7052 4324 7058 4326
rect 7114 4324 7138 4326
rect 7194 4324 7218 4326
rect 7274 4324 7298 4326
rect 7354 4324 7360 4326
rect 7052 4304 7360 4324
rect 7484 4146 7512 4558
rect 9140 4486 9168 5578
rect 9324 4622 9352 5714
rect 9404 5704 9456 5710
rect 9456 5664 9536 5692
rect 9404 5646 9456 5652
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5302 9444 5510
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9508 5166 9536 5664
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9600 5148 9628 6938
rect 9968 6798 9996 7482
rect 10104 7100 10412 7120
rect 10104 7098 10110 7100
rect 10166 7098 10190 7100
rect 10246 7098 10270 7100
rect 10326 7098 10350 7100
rect 10406 7098 10412 7100
rect 10166 7046 10168 7098
rect 10348 7046 10350 7098
rect 10104 7044 10110 7046
rect 10166 7044 10190 7046
rect 10246 7044 10270 7046
rect 10326 7044 10350 7046
rect 10406 7044 10412 7046
rect 10104 7024 10412 7044
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10104 6012 10412 6032
rect 10104 6010 10110 6012
rect 10166 6010 10190 6012
rect 10246 6010 10270 6012
rect 10326 6010 10350 6012
rect 10406 6010 10412 6012
rect 10166 5958 10168 6010
rect 10348 5958 10350 6010
rect 10104 5956 10110 5958
rect 10166 5956 10190 5958
rect 10246 5956 10270 5958
rect 10326 5956 10350 5958
rect 10406 5956 10412 5958
rect 10104 5936 10412 5956
rect 10888 5710 10916 7686
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 9772 5160 9824 5166
rect 9600 5120 9772 5148
rect 9508 4826 9536 5102
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9600 4690 9628 5120
rect 9772 5102 9824 5108
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3126 6868 3334
rect 7052 3292 7360 3312
rect 7052 3290 7058 3292
rect 7114 3290 7138 3292
rect 7194 3290 7218 3292
rect 7274 3290 7298 3292
rect 7354 3290 7360 3292
rect 7114 3238 7116 3290
rect 7296 3238 7298 3290
rect 7052 3236 7058 3238
rect 7114 3236 7138 3238
rect 7194 3236 7218 3238
rect 7274 3236 7298 3238
rect 7354 3236 7360 3238
rect 7052 3216 7360 3236
rect 7392 3126 7420 3878
rect 7484 3602 7512 3878
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7852 3534 7880 4422
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8036 3534 8064 4014
rect 8128 3602 8156 4082
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8036 3176 8064 3470
rect 8116 3188 8168 3194
rect 8036 3148 8116 3176
rect 8116 3130 8168 3136
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 9600 3058 9628 4626
rect 9968 3602 9996 4966
rect 10104 4924 10412 4944
rect 10104 4922 10110 4924
rect 10166 4922 10190 4924
rect 10246 4922 10270 4924
rect 10326 4922 10350 4924
rect 10406 4922 10412 4924
rect 10166 4870 10168 4922
rect 10348 4870 10350 4922
rect 10104 4868 10110 4870
rect 10166 4868 10190 4870
rect 10246 4868 10270 4870
rect 10326 4868 10350 4870
rect 10406 4868 10412 4870
rect 10104 4848 10412 4868
rect 10888 4690 10916 5646
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10104 3836 10412 3856
rect 10104 3834 10110 3836
rect 10166 3834 10190 3836
rect 10246 3834 10270 3836
rect 10326 3834 10350 3836
rect 10406 3834 10412 3836
rect 10166 3782 10168 3834
rect 10348 3782 10350 3834
rect 10104 3780 10110 3782
rect 10166 3780 10190 3782
rect 10246 3780 10270 3782
rect 10326 3780 10350 3782
rect 10406 3780 10412 3782
rect 10104 3760 10412 3780
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 3194 9812 3402
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 10980 3040 11008 7278
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 5914 12388 6190
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12452 5778 12480 6802
rect 12544 6746 12572 9318
rect 12636 7954 12664 10474
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12728 7410 12756 8366
rect 12820 8090 12848 8502
rect 12912 8294 12940 10066
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12912 7954 12940 8230
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 13004 7886 13032 11086
rect 13155 10908 13463 10928
rect 13155 10906 13161 10908
rect 13217 10906 13241 10908
rect 13297 10906 13321 10908
rect 13377 10906 13401 10908
rect 13457 10906 13463 10908
rect 13217 10854 13219 10906
rect 13399 10854 13401 10906
rect 13155 10852 13161 10854
rect 13217 10852 13241 10854
rect 13297 10852 13321 10854
rect 13377 10852 13401 10854
rect 13457 10852 13463 10854
rect 13155 10832 13463 10852
rect 13556 10742 13584 11086
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13155 9820 13463 9840
rect 13155 9818 13161 9820
rect 13217 9818 13241 9820
rect 13297 9818 13321 9820
rect 13377 9818 13401 9820
rect 13457 9818 13463 9820
rect 13217 9766 13219 9818
rect 13399 9766 13401 9818
rect 13155 9764 13161 9766
rect 13217 9764 13241 9766
rect 13297 9764 13321 9766
rect 13377 9764 13401 9766
rect 13457 9764 13463 9766
rect 13155 9744 13463 9764
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13155 8732 13463 8752
rect 13155 8730 13161 8732
rect 13217 8730 13241 8732
rect 13297 8730 13321 8732
rect 13377 8730 13401 8732
rect 13457 8730 13463 8732
rect 13217 8678 13219 8730
rect 13399 8678 13401 8730
rect 13155 8676 13161 8678
rect 13217 8676 13241 8678
rect 13297 8676 13321 8678
rect 13377 8676 13401 8678
rect 13457 8676 13463 8678
rect 13155 8656 13463 8676
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 6866 12756 7346
rect 13004 7274 13032 7822
rect 13155 7644 13463 7664
rect 13155 7642 13161 7644
rect 13217 7642 13241 7644
rect 13297 7642 13321 7644
rect 13377 7642 13401 7644
rect 13457 7642 13463 7644
rect 13217 7590 13219 7642
rect 13399 7590 13401 7642
rect 13155 7588 13161 7590
rect 13217 7588 13241 7590
rect 13297 7588 13321 7590
rect 13377 7588 13401 7590
rect 13457 7588 13463 7590
rect 13155 7568 13463 7588
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12544 6718 12756 6746
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5370 11100 5646
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11072 4622 11100 5306
rect 12452 5166 12480 5714
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 12544 4146 12572 6054
rect 12728 5846 12756 6718
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12728 5710 12756 5782
rect 12820 5778 12848 7142
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12544 3602 12572 4082
rect 12636 4026 12664 4558
rect 12728 4214 12756 5034
rect 12912 4826 12940 6258
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12636 3998 12756 4026
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12544 3058 12572 3538
rect 12728 3466 12756 3998
rect 13004 3738 13032 7210
rect 13096 6798 13124 7346
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6458 13124 6734
rect 13155 6556 13463 6576
rect 13155 6554 13161 6556
rect 13217 6554 13241 6556
rect 13297 6554 13321 6556
rect 13377 6554 13401 6556
rect 13457 6554 13463 6556
rect 13217 6502 13219 6554
rect 13399 6502 13401 6554
rect 13155 6500 13161 6502
rect 13217 6500 13241 6502
rect 13297 6500 13321 6502
rect 13377 6500 13401 6502
rect 13457 6500 13463 6502
rect 13155 6480 13463 6500
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13740 6322 13768 8298
rect 13832 7410 13860 8842
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13155 5468 13463 5488
rect 13155 5466 13161 5468
rect 13217 5466 13241 5468
rect 13297 5466 13321 5468
rect 13377 5466 13401 5468
rect 13457 5466 13463 5468
rect 13217 5414 13219 5466
rect 13399 5414 13401 5466
rect 13155 5412 13161 5414
rect 13217 5412 13241 5414
rect 13297 5412 13321 5414
rect 13377 5412 13401 5414
rect 13457 5412 13463 5414
rect 13155 5392 13463 5412
rect 13556 5234 13584 5510
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13924 4690 13952 12406
rect 14016 12238 14044 12854
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14016 11762 14044 12174
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14016 9994 14044 11698
rect 14200 11626 14228 13874
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14752 12850 14780 13330
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12434 14412 12582
rect 14384 12406 14504 12434
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11218 14136 11494
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14108 10742 14136 11154
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 14016 9654 14044 9930
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14108 9382 14136 10406
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 8362 14136 9318
rect 14200 8974 14228 11562
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14292 8566 14320 8774
rect 14384 8634 14412 8774
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14108 7954 14136 8298
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14476 6746 14504 12406
rect 14752 12306 14780 12786
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14752 11898 14780 12242
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 11762 14872 13806
rect 15120 13190 15148 13874
rect 15396 13530 15424 14282
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12850 15148 13126
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14752 7546 14780 9590
rect 14844 9178 14872 11698
rect 15580 11234 15608 19790
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15672 18834 15700 19110
rect 15856 18902 15884 19110
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15856 18766 15884 18838
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15764 16522 15792 16934
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15856 15586 15884 18090
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15948 16250 15976 17614
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15764 15558 15884 15586
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15672 12986 15700 15030
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15672 12306 15700 12922
rect 15764 12434 15792 15558
rect 16040 15502 16068 18906
rect 16132 18834 16160 21950
rect 16394 21861 16450 21950
rect 17038 21861 17094 22661
rect 17682 21861 17738 22661
rect 18234 21861 18290 22661
rect 18878 21861 18934 22661
rect 19522 21861 19578 22661
rect 20166 21861 20222 22661
rect 16206 20156 16514 20176
rect 16206 20154 16212 20156
rect 16268 20154 16292 20156
rect 16348 20154 16372 20156
rect 16428 20154 16452 20156
rect 16508 20154 16514 20156
rect 16268 20102 16270 20154
rect 16450 20102 16452 20154
rect 16206 20100 16212 20102
rect 16268 20100 16292 20102
rect 16348 20100 16372 20102
rect 16428 20100 16452 20102
rect 16508 20100 16514 20102
rect 16206 20080 16514 20100
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16206 19068 16514 19088
rect 16206 19066 16212 19068
rect 16268 19066 16292 19068
rect 16348 19066 16372 19068
rect 16428 19066 16452 19068
rect 16508 19066 16514 19068
rect 16268 19014 16270 19066
rect 16450 19014 16452 19066
rect 16206 19012 16212 19014
rect 16268 19012 16292 19014
rect 16348 19012 16372 19014
rect 16428 19012 16452 19014
rect 16508 19012 16514 19014
rect 16206 18992 16514 19012
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16132 17610 16160 18158
rect 16206 17980 16514 18000
rect 16206 17978 16212 17980
rect 16268 17978 16292 17980
rect 16348 17978 16372 17980
rect 16428 17978 16452 17980
rect 16508 17978 16514 17980
rect 16268 17926 16270 17978
rect 16450 17926 16452 17978
rect 16206 17924 16212 17926
rect 16268 17924 16292 17926
rect 16348 17924 16372 17926
rect 16428 17924 16452 17926
rect 16508 17924 16514 17926
rect 16206 17904 16514 17924
rect 16592 17882 16620 18294
rect 16684 18290 16712 19450
rect 17052 18834 17080 21861
rect 17696 19922 17724 21861
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 16592 17338 16620 17614
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16206 16892 16514 16912
rect 16206 16890 16212 16892
rect 16268 16890 16292 16892
rect 16348 16890 16372 16892
rect 16428 16890 16452 16892
rect 16508 16890 16514 16892
rect 16268 16838 16270 16890
rect 16450 16838 16452 16890
rect 16206 16836 16212 16838
rect 16268 16836 16292 16838
rect 16348 16836 16372 16838
rect 16428 16836 16452 16838
rect 16508 16836 16514 16838
rect 16206 16816 16514 16836
rect 16684 16658 16712 18226
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16960 17882 16988 18158
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16206 15804 16514 15824
rect 16206 15802 16212 15804
rect 16268 15802 16292 15804
rect 16348 15802 16372 15804
rect 16428 15802 16452 15804
rect 16508 15802 16514 15804
rect 16268 15750 16270 15802
rect 16450 15750 16452 15802
rect 16206 15748 16212 15750
rect 16268 15748 16292 15750
rect 16348 15748 16372 15750
rect 16428 15748 16452 15750
rect 16508 15748 16514 15750
rect 16206 15728 16514 15748
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15856 15026 15884 15438
rect 16592 15366 16620 16050
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15856 14618 15884 14962
rect 16206 14716 16514 14736
rect 16206 14714 16212 14716
rect 16268 14714 16292 14716
rect 16348 14714 16372 14716
rect 16428 14714 16452 14716
rect 16508 14714 16514 14716
rect 16268 14662 16270 14714
rect 16450 14662 16452 14714
rect 16206 14660 16212 14662
rect 16268 14660 16292 14662
rect 16348 14660 16372 14662
rect 16428 14660 16452 14662
rect 16508 14660 16514 14662
rect 16206 14640 16514 14660
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 16592 14074 16620 15098
rect 16684 15026 16712 16594
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16684 14482 16712 14962
rect 16776 14482 16804 15302
rect 16868 14550 16896 15914
rect 16960 15502 16988 17138
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16960 15162 16988 15438
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14618 16988 14894
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16206 13628 16514 13648
rect 16206 13626 16212 13628
rect 16268 13626 16292 13628
rect 16348 13626 16372 13628
rect 16428 13626 16452 13628
rect 16508 13626 16514 13628
rect 16268 13574 16270 13626
rect 16450 13574 16452 13626
rect 16206 13572 16212 13574
rect 16268 13572 16292 13574
rect 16348 13572 16372 13574
rect 16428 13572 16452 13574
rect 16508 13572 16514 13574
rect 16206 13552 16514 13572
rect 16684 13394 16712 14418
rect 16868 14414 16896 14486
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 17052 13938 17080 18022
rect 17144 16130 17172 19790
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17236 16250 17264 16458
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17144 16102 17264 16130
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17144 14482 17172 15370
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16040 12434 16068 13330
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 12986 16160 13262
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16206 12540 16514 12560
rect 16206 12538 16212 12540
rect 16268 12538 16292 12540
rect 16348 12538 16372 12540
rect 16428 12538 16452 12540
rect 16508 12538 16514 12540
rect 16268 12486 16270 12538
rect 16450 12486 16452 12538
rect 16206 12484 16212 12486
rect 16268 12484 16292 12486
rect 16348 12484 16372 12486
rect 16428 12484 16452 12486
rect 16508 12484 16514 12486
rect 16206 12464 16514 12484
rect 15764 12406 15884 12434
rect 16040 12406 16252 12434
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15856 12186 15884 12406
rect 16224 12238 16252 12406
rect 16212 12232 16264 12238
rect 15856 12158 16068 12186
rect 16212 12174 16264 12180
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15842 11248 15898 11257
rect 15580 11206 15792 11234
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10674 15240 10950
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9518 14964 9862
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 15120 8974 15148 9454
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15212 8498 15240 10610
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10130 15424 10542
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15488 10130 15516 10474
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15396 9178 15424 10066
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15580 8974 15608 11086
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15672 9722 15700 9998
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15396 7954 15424 8570
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7546 15516 7822
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15028 7206 15056 7346
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6798 15056 7142
rect 14292 6718 14504 6746
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14292 5166 14320 6718
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 14936 6390 14964 6598
rect 15672 6458 15700 6598
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15764 6390 15792 11206
rect 15842 11183 15898 11192
rect 15856 11082 15884 11183
rect 15948 11082 15976 12038
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 16040 10146 16068 12158
rect 16224 11694 16252 12174
rect 16776 11762 16804 12718
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16206 11452 16514 11472
rect 16206 11450 16212 11452
rect 16268 11450 16292 11452
rect 16348 11450 16372 11452
rect 16428 11450 16452 11452
rect 16508 11450 16514 11452
rect 16268 11398 16270 11450
rect 16450 11398 16452 11450
rect 16206 11396 16212 11398
rect 16268 11396 16292 11398
rect 16348 11396 16372 11398
rect 16428 11396 16452 11398
rect 16508 11396 16514 11398
rect 16206 11376 16514 11396
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16592 10606 16620 11154
rect 16684 11082 16712 11494
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16206 10364 16514 10384
rect 16206 10362 16212 10364
rect 16268 10362 16292 10364
rect 16348 10362 16372 10364
rect 16428 10362 16452 10364
rect 16508 10362 16514 10364
rect 16268 10310 16270 10362
rect 16450 10310 16452 10362
rect 16206 10308 16212 10310
rect 16268 10308 16292 10310
rect 16348 10308 16372 10310
rect 16428 10308 16452 10310
rect 16508 10308 16514 10310
rect 16206 10288 16514 10308
rect 15948 10118 16068 10146
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15856 9110 15884 9522
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15856 8090 15884 9046
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5710 15608 6190
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15948 5574 15976 10118
rect 16776 10062 16804 11698
rect 17236 10606 17264 16102
rect 17328 15162 17356 17546
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17512 15502 17540 16050
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17328 14414 17356 15098
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17328 11014 17356 12786
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 16040 8906 16068 9930
rect 16206 9276 16514 9296
rect 16206 9274 16212 9276
rect 16268 9274 16292 9276
rect 16348 9274 16372 9276
rect 16428 9274 16452 9276
rect 16508 9274 16514 9276
rect 16268 9222 16270 9274
rect 16450 9222 16452 9274
rect 16206 9220 16212 9222
rect 16268 9220 16292 9222
rect 16348 9220 16372 9222
rect 16428 9220 16452 9222
rect 16508 9220 16514 9222
rect 16206 9200 16514 9220
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 16040 6866 16068 8842
rect 16592 8498 16620 8978
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16206 8188 16514 8208
rect 16206 8186 16212 8188
rect 16268 8186 16292 8188
rect 16348 8186 16372 8188
rect 16428 8186 16452 8188
rect 16508 8186 16514 8188
rect 16268 8134 16270 8186
rect 16450 8134 16452 8186
rect 16206 8132 16212 8134
rect 16268 8132 16292 8134
rect 16348 8132 16372 8134
rect 16428 8132 16452 8134
rect 16508 8132 16514 8134
rect 16206 8112 16514 8132
rect 16776 7342 16804 9998
rect 16868 9518 16896 10542
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 16868 8820 16896 9454
rect 17144 9178 17172 9454
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 16868 8792 16988 8820
rect 16960 8294 16988 8792
rect 17144 8430 17172 8910
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16960 7342 16988 8230
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 16206 7100 16514 7120
rect 16206 7098 16212 7100
rect 16268 7098 16292 7100
rect 16348 7098 16372 7100
rect 16428 7098 16452 7100
rect 16508 7098 16514 7100
rect 16268 7046 16270 7098
rect 16450 7046 16452 7098
rect 16206 7044 16212 7046
rect 16268 7044 16292 7046
rect 16348 7044 16372 7046
rect 16428 7044 16452 7046
rect 16508 7044 16514 7046
rect 16206 7024 16514 7044
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 14292 4622 14320 5102
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13155 4380 13463 4400
rect 13155 4378 13161 4380
rect 13217 4378 13241 4380
rect 13297 4378 13321 4380
rect 13377 4378 13401 4380
rect 13457 4378 13463 4380
rect 13217 4326 13219 4378
rect 13399 4326 13401 4378
rect 13155 4324 13161 4326
rect 13217 4324 13241 4326
rect 13297 4324 13321 4326
rect 13377 4324 13401 4326
rect 13457 4324 13463 4326
rect 13155 4304 13463 4324
rect 13556 4214 13584 4422
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 14476 4078 14504 4558
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 11060 3052 11112 3058
rect 10980 3012 11060 3040
rect 10980 2774 11008 3012
rect 11060 2994 11112 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12728 2990 12756 3402
rect 13155 3292 13463 3312
rect 13155 3290 13161 3292
rect 13217 3290 13241 3292
rect 13297 3290 13321 3292
rect 13377 3290 13401 3292
rect 13457 3290 13463 3292
rect 13217 3238 13219 3290
rect 13399 3238 13401 3290
rect 13155 3236 13161 3238
rect 13217 3236 13241 3238
rect 13297 3236 13321 3238
rect 13377 3236 13401 3238
rect 13457 3236 13463 3238
rect 13155 3216 13463 3236
rect 14568 3194 14596 3878
rect 14752 3534 14780 5102
rect 14936 4282 14964 5170
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14936 3602 14964 4218
rect 15028 4146 15056 4626
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 15028 3738 15056 4082
rect 15212 4078 15240 4490
rect 15304 4146 15332 4966
rect 16040 4554 16068 6802
rect 16132 5914 16160 6870
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6458 16712 6734
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16206 6012 16514 6032
rect 16206 6010 16212 6012
rect 16268 6010 16292 6012
rect 16348 6010 16372 6012
rect 16428 6010 16452 6012
rect 16508 6010 16514 6012
rect 16268 5958 16270 6010
rect 16450 5958 16452 6010
rect 16206 5956 16212 5958
rect 16268 5956 16292 5958
rect 16348 5956 16372 5958
rect 16428 5956 16452 5958
rect 16508 5956 16514 5958
rect 16206 5936 16514 5956
rect 16868 5914 16896 6258
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16960 5710 16988 7278
rect 17236 6934 17264 7278
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17328 6798 17356 10950
rect 17604 9042 17632 18702
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17696 15706 17724 16458
rect 17972 16250 18000 19382
rect 18064 18442 18092 19858
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18156 18714 18184 19790
rect 18248 19786 18276 21861
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18524 19446 18552 19654
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18328 18760 18380 18766
rect 18156 18686 18276 18714
rect 18328 18702 18380 18708
rect 18064 18414 18184 18442
rect 18156 17762 18184 18414
rect 18248 17814 18276 18686
rect 18064 17746 18184 17762
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18052 17740 18184 17746
rect 18104 17734 18184 17740
rect 18052 17682 18104 17688
rect 18064 17066 18092 17682
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 15094 18000 15302
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17972 12850 18000 14010
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11354 17908 12174
rect 17972 12170 18000 12786
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 18156 11830 18184 17614
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18248 16794 18276 17070
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18248 14482 18276 15438
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17972 11218 18000 11698
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 18064 11150 18092 11562
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18064 10810 18092 11086
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17972 10266 18000 10678
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9654 18184 9862
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18156 7546 18184 7822
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18156 7290 18184 7482
rect 18248 7478 18276 7686
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18156 7262 18276 7290
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17696 6322 17724 6734
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16206 4924 16514 4944
rect 16206 4922 16212 4924
rect 16268 4922 16292 4924
rect 16348 4922 16372 4924
rect 16428 4922 16452 4924
rect 16508 4922 16514 4924
rect 16268 4870 16270 4922
rect 16450 4870 16452 4922
rect 16206 4868 16212 4870
rect 16268 4868 16292 4870
rect 16348 4868 16372 4870
rect 16428 4868 16452 4870
rect 16508 4868 16514 4870
rect 16206 4848 16514 4868
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3194 14780 3470
rect 15764 3466 15792 4422
rect 16592 4078 16620 5646
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17236 5370 17264 5578
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17420 5234 17448 6054
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17328 4622 17356 5102
rect 17512 4758 17540 6258
rect 18248 5234 18276 7262
rect 18340 6798 18368 18702
rect 18892 18426 18920 21861
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18432 17202 18460 18022
rect 19536 17746 19564 21861
rect 20180 19990 20208 21861
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18432 15162 18460 15438
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18432 14414 18460 15098
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18708 13530 18736 14418
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18524 12986 18552 13194
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 9042 18552 9318
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18524 8498 18552 8978
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18708 8430 18736 8910
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18708 7546 18736 8366
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18340 5370 18368 5646
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 17500 4752 17552 4758
rect 17500 4694 17552 4700
rect 18248 4622 18276 5170
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16960 4214 16988 4422
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16206 3836 16514 3856
rect 16206 3834 16212 3836
rect 16268 3834 16292 3836
rect 16348 3834 16372 3836
rect 16428 3834 16452 3836
rect 16508 3834 16514 3836
rect 16268 3782 16270 3834
rect 16450 3782 16452 3834
rect 16206 3780 16212 3782
rect 16268 3780 16292 3782
rect 16348 3780 16372 3782
rect 16428 3780 16452 3782
rect 16508 3780 16514 3782
rect 16206 3760 16514 3780
rect 16592 3618 16620 4014
rect 17328 3738 17356 4558
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 16500 3602 16620 3618
rect 16488 3596 16620 3602
rect 16540 3590 16620 3596
rect 16488 3538 16540 3544
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16224 3194 16252 3402
rect 17604 3194 17632 4558
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18248 4214 18276 4422
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 4001 2748 4309 2768
rect 4001 2746 4007 2748
rect 4063 2746 4087 2748
rect 4143 2746 4167 2748
rect 4223 2746 4247 2748
rect 4303 2746 4309 2748
rect 4063 2694 4065 2746
rect 4245 2694 4247 2746
rect 4001 2692 4007 2694
rect 4063 2692 4087 2694
rect 4143 2692 4167 2694
rect 4223 2692 4247 2694
rect 4303 2692 4309 2694
rect 4001 2672 4309 2692
rect 10104 2748 10412 2768
rect 10104 2746 10110 2748
rect 10166 2746 10190 2748
rect 10246 2746 10270 2748
rect 10326 2746 10350 2748
rect 10406 2746 10412 2748
rect 10166 2694 10168 2746
rect 10348 2694 10350 2746
rect 10104 2692 10110 2694
rect 10166 2692 10190 2694
rect 10246 2692 10270 2694
rect 10326 2692 10350 2694
rect 10406 2692 10412 2694
rect 10104 2672 10412 2692
rect 10612 2746 11008 2774
rect 10612 2582 10640 2746
rect 14292 2650 14320 3062
rect 17788 3058 17816 3606
rect 18064 3534 18092 3878
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18064 3058 18092 3470
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 14568 2446 14596 2994
rect 16206 2748 16514 2768
rect 16206 2746 16212 2748
rect 16268 2746 16292 2748
rect 16348 2746 16372 2748
rect 16428 2746 16452 2748
rect 16508 2746 16514 2748
rect 16268 2694 16270 2746
rect 16450 2694 16452 2746
rect 16206 2692 16212 2694
rect 16268 2692 16292 2694
rect 16348 2692 16372 2694
rect 16428 2692 16452 2694
rect 16508 2692 16514 2694
rect 16206 2672 16514 2692
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 7052 2204 7360 2224
rect 7052 2202 7058 2204
rect 7114 2202 7138 2204
rect 7194 2202 7218 2204
rect 7274 2202 7298 2204
rect 7354 2202 7360 2204
rect 7114 2150 7116 2202
rect 7296 2150 7298 2202
rect 7052 2148 7058 2150
rect 7114 2148 7138 2150
rect 7194 2148 7218 2150
rect 7274 2148 7298 2150
rect 7354 2148 7360 2150
rect 7052 2128 7360 2148
rect 10244 800 10272 2314
rect 13155 2204 13463 2224
rect 13155 2202 13161 2204
rect 13217 2202 13241 2204
rect 13297 2202 13321 2204
rect 13377 2202 13401 2204
rect 13457 2202 13463 2204
rect 13217 2150 13219 2202
rect 13399 2150 13401 2202
rect 13155 2148 13161 2150
rect 13217 2148 13241 2150
rect 13297 2148 13321 2150
rect 13377 2148 13401 2150
rect 13457 2148 13463 2150
rect 13155 2128 13463 2148
rect 10230 0 10286 800
<< via2 >>
rect 1582 11328 1638 11384
rect 4007 20154 4063 20156
rect 4087 20154 4143 20156
rect 4167 20154 4223 20156
rect 4247 20154 4303 20156
rect 4007 20102 4053 20154
rect 4053 20102 4063 20154
rect 4087 20102 4117 20154
rect 4117 20102 4129 20154
rect 4129 20102 4143 20154
rect 4167 20102 4181 20154
rect 4181 20102 4193 20154
rect 4193 20102 4223 20154
rect 4247 20102 4257 20154
rect 4257 20102 4303 20154
rect 4007 20100 4063 20102
rect 4087 20100 4143 20102
rect 4167 20100 4223 20102
rect 4247 20100 4303 20102
rect 4007 19066 4063 19068
rect 4087 19066 4143 19068
rect 4167 19066 4223 19068
rect 4247 19066 4303 19068
rect 4007 19014 4053 19066
rect 4053 19014 4063 19066
rect 4087 19014 4117 19066
rect 4117 19014 4129 19066
rect 4129 19014 4143 19066
rect 4167 19014 4181 19066
rect 4181 19014 4193 19066
rect 4193 19014 4223 19066
rect 4247 19014 4257 19066
rect 4257 19014 4303 19066
rect 4007 19012 4063 19014
rect 4087 19012 4143 19014
rect 4167 19012 4223 19014
rect 4247 19012 4303 19014
rect 4007 17978 4063 17980
rect 4087 17978 4143 17980
rect 4167 17978 4223 17980
rect 4247 17978 4303 17980
rect 4007 17926 4053 17978
rect 4053 17926 4063 17978
rect 4087 17926 4117 17978
rect 4117 17926 4129 17978
rect 4129 17926 4143 17978
rect 4167 17926 4181 17978
rect 4181 17926 4193 17978
rect 4193 17926 4223 17978
rect 4247 17926 4257 17978
rect 4257 17926 4303 17978
rect 4007 17924 4063 17926
rect 4087 17924 4143 17926
rect 4167 17924 4223 17926
rect 4247 17924 4303 17926
rect 4007 16890 4063 16892
rect 4087 16890 4143 16892
rect 4167 16890 4223 16892
rect 4247 16890 4303 16892
rect 4007 16838 4053 16890
rect 4053 16838 4063 16890
rect 4087 16838 4117 16890
rect 4117 16838 4129 16890
rect 4129 16838 4143 16890
rect 4167 16838 4181 16890
rect 4181 16838 4193 16890
rect 4193 16838 4223 16890
rect 4247 16838 4257 16890
rect 4257 16838 4303 16890
rect 4007 16836 4063 16838
rect 4087 16836 4143 16838
rect 4167 16836 4223 16838
rect 4247 16836 4303 16838
rect 4007 15802 4063 15804
rect 4087 15802 4143 15804
rect 4167 15802 4223 15804
rect 4247 15802 4303 15804
rect 4007 15750 4053 15802
rect 4053 15750 4063 15802
rect 4087 15750 4117 15802
rect 4117 15750 4129 15802
rect 4129 15750 4143 15802
rect 4167 15750 4181 15802
rect 4181 15750 4193 15802
rect 4193 15750 4223 15802
rect 4247 15750 4257 15802
rect 4257 15750 4303 15802
rect 4007 15748 4063 15750
rect 4087 15748 4143 15750
rect 4167 15748 4223 15750
rect 4247 15748 4303 15750
rect 4007 14714 4063 14716
rect 4087 14714 4143 14716
rect 4167 14714 4223 14716
rect 4247 14714 4303 14716
rect 4007 14662 4053 14714
rect 4053 14662 4063 14714
rect 4087 14662 4117 14714
rect 4117 14662 4129 14714
rect 4129 14662 4143 14714
rect 4167 14662 4181 14714
rect 4181 14662 4193 14714
rect 4193 14662 4223 14714
rect 4247 14662 4257 14714
rect 4257 14662 4303 14714
rect 4007 14660 4063 14662
rect 4087 14660 4143 14662
rect 4167 14660 4223 14662
rect 4247 14660 4303 14662
rect 4007 13626 4063 13628
rect 4087 13626 4143 13628
rect 4167 13626 4223 13628
rect 4247 13626 4303 13628
rect 4007 13574 4053 13626
rect 4053 13574 4063 13626
rect 4087 13574 4117 13626
rect 4117 13574 4129 13626
rect 4129 13574 4143 13626
rect 4167 13574 4181 13626
rect 4181 13574 4193 13626
rect 4193 13574 4223 13626
rect 4247 13574 4257 13626
rect 4257 13574 4303 13626
rect 4007 13572 4063 13574
rect 4087 13572 4143 13574
rect 4167 13572 4223 13574
rect 4247 13572 4303 13574
rect 4007 12538 4063 12540
rect 4087 12538 4143 12540
rect 4167 12538 4223 12540
rect 4247 12538 4303 12540
rect 4007 12486 4053 12538
rect 4053 12486 4063 12538
rect 4087 12486 4117 12538
rect 4117 12486 4129 12538
rect 4129 12486 4143 12538
rect 4167 12486 4181 12538
rect 4181 12486 4193 12538
rect 4193 12486 4223 12538
rect 4247 12486 4257 12538
rect 4257 12486 4303 12538
rect 4007 12484 4063 12486
rect 4087 12484 4143 12486
rect 4167 12484 4223 12486
rect 4247 12484 4303 12486
rect 4007 11450 4063 11452
rect 4087 11450 4143 11452
rect 4167 11450 4223 11452
rect 4247 11450 4303 11452
rect 4007 11398 4053 11450
rect 4053 11398 4063 11450
rect 4087 11398 4117 11450
rect 4117 11398 4129 11450
rect 4129 11398 4143 11450
rect 4167 11398 4181 11450
rect 4181 11398 4193 11450
rect 4193 11398 4223 11450
rect 4247 11398 4257 11450
rect 4257 11398 4303 11450
rect 4007 11396 4063 11398
rect 4087 11396 4143 11398
rect 4167 11396 4223 11398
rect 4247 11396 4303 11398
rect 4007 10362 4063 10364
rect 4087 10362 4143 10364
rect 4167 10362 4223 10364
rect 4247 10362 4303 10364
rect 4007 10310 4053 10362
rect 4053 10310 4063 10362
rect 4087 10310 4117 10362
rect 4117 10310 4129 10362
rect 4129 10310 4143 10362
rect 4167 10310 4181 10362
rect 4181 10310 4193 10362
rect 4193 10310 4223 10362
rect 4247 10310 4257 10362
rect 4257 10310 4303 10362
rect 4007 10308 4063 10310
rect 4087 10308 4143 10310
rect 4167 10308 4223 10310
rect 4247 10308 4303 10310
rect 4007 9274 4063 9276
rect 4087 9274 4143 9276
rect 4167 9274 4223 9276
rect 4247 9274 4303 9276
rect 4007 9222 4053 9274
rect 4053 9222 4063 9274
rect 4087 9222 4117 9274
rect 4117 9222 4129 9274
rect 4129 9222 4143 9274
rect 4167 9222 4181 9274
rect 4181 9222 4193 9274
rect 4193 9222 4223 9274
rect 4247 9222 4257 9274
rect 4257 9222 4303 9274
rect 4007 9220 4063 9222
rect 4087 9220 4143 9222
rect 4167 9220 4223 9222
rect 4247 9220 4303 9222
rect 4007 8186 4063 8188
rect 4087 8186 4143 8188
rect 4167 8186 4223 8188
rect 4247 8186 4303 8188
rect 4007 8134 4053 8186
rect 4053 8134 4063 8186
rect 4087 8134 4117 8186
rect 4117 8134 4129 8186
rect 4129 8134 4143 8186
rect 4167 8134 4181 8186
rect 4181 8134 4193 8186
rect 4193 8134 4223 8186
rect 4247 8134 4257 8186
rect 4257 8134 4303 8186
rect 4007 8132 4063 8134
rect 4087 8132 4143 8134
rect 4167 8132 4223 8134
rect 4247 8132 4303 8134
rect 4007 7098 4063 7100
rect 4087 7098 4143 7100
rect 4167 7098 4223 7100
rect 4247 7098 4303 7100
rect 4007 7046 4053 7098
rect 4053 7046 4063 7098
rect 4087 7046 4117 7098
rect 4117 7046 4129 7098
rect 4129 7046 4143 7098
rect 4167 7046 4181 7098
rect 4181 7046 4193 7098
rect 4193 7046 4223 7098
rect 4247 7046 4257 7098
rect 4257 7046 4303 7098
rect 4007 7044 4063 7046
rect 4087 7044 4143 7046
rect 4167 7044 4223 7046
rect 4247 7044 4303 7046
rect 7058 19610 7114 19612
rect 7138 19610 7194 19612
rect 7218 19610 7274 19612
rect 7298 19610 7354 19612
rect 7058 19558 7104 19610
rect 7104 19558 7114 19610
rect 7138 19558 7168 19610
rect 7168 19558 7180 19610
rect 7180 19558 7194 19610
rect 7218 19558 7232 19610
rect 7232 19558 7244 19610
rect 7244 19558 7274 19610
rect 7298 19558 7308 19610
rect 7308 19558 7354 19610
rect 7058 19556 7114 19558
rect 7138 19556 7194 19558
rect 7218 19556 7274 19558
rect 7298 19556 7354 19558
rect 7058 18522 7114 18524
rect 7138 18522 7194 18524
rect 7218 18522 7274 18524
rect 7298 18522 7354 18524
rect 7058 18470 7104 18522
rect 7104 18470 7114 18522
rect 7138 18470 7168 18522
rect 7168 18470 7180 18522
rect 7180 18470 7194 18522
rect 7218 18470 7232 18522
rect 7232 18470 7244 18522
rect 7244 18470 7274 18522
rect 7298 18470 7308 18522
rect 7308 18470 7354 18522
rect 7058 18468 7114 18470
rect 7138 18468 7194 18470
rect 7218 18468 7274 18470
rect 7298 18468 7354 18470
rect 7058 17434 7114 17436
rect 7138 17434 7194 17436
rect 7218 17434 7274 17436
rect 7298 17434 7354 17436
rect 7058 17382 7104 17434
rect 7104 17382 7114 17434
rect 7138 17382 7168 17434
rect 7168 17382 7180 17434
rect 7180 17382 7194 17434
rect 7218 17382 7232 17434
rect 7232 17382 7244 17434
rect 7244 17382 7274 17434
rect 7298 17382 7308 17434
rect 7308 17382 7354 17434
rect 7058 17380 7114 17382
rect 7138 17380 7194 17382
rect 7218 17380 7274 17382
rect 7298 17380 7354 17382
rect 7058 16346 7114 16348
rect 7138 16346 7194 16348
rect 7218 16346 7274 16348
rect 7298 16346 7354 16348
rect 7058 16294 7104 16346
rect 7104 16294 7114 16346
rect 7138 16294 7168 16346
rect 7168 16294 7180 16346
rect 7180 16294 7194 16346
rect 7218 16294 7232 16346
rect 7232 16294 7244 16346
rect 7244 16294 7274 16346
rect 7298 16294 7308 16346
rect 7308 16294 7354 16346
rect 7058 16292 7114 16294
rect 7138 16292 7194 16294
rect 7218 16292 7274 16294
rect 7298 16292 7354 16294
rect 7058 15258 7114 15260
rect 7138 15258 7194 15260
rect 7218 15258 7274 15260
rect 7298 15258 7354 15260
rect 7058 15206 7104 15258
rect 7104 15206 7114 15258
rect 7138 15206 7168 15258
rect 7168 15206 7180 15258
rect 7180 15206 7194 15258
rect 7218 15206 7232 15258
rect 7232 15206 7244 15258
rect 7244 15206 7274 15258
rect 7298 15206 7308 15258
rect 7308 15206 7354 15258
rect 7058 15204 7114 15206
rect 7138 15204 7194 15206
rect 7218 15204 7274 15206
rect 7298 15204 7354 15206
rect 4007 6010 4063 6012
rect 4087 6010 4143 6012
rect 4167 6010 4223 6012
rect 4247 6010 4303 6012
rect 4007 5958 4053 6010
rect 4053 5958 4063 6010
rect 4087 5958 4117 6010
rect 4117 5958 4129 6010
rect 4129 5958 4143 6010
rect 4167 5958 4181 6010
rect 4181 5958 4193 6010
rect 4193 5958 4223 6010
rect 4247 5958 4257 6010
rect 4257 5958 4303 6010
rect 4007 5956 4063 5958
rect 4087 5956 4143 5958
rect 4167 5956 4223 5958
rect 4247 5956 4303 5958
rect 7058 14170 7114 14172
rect 7138 14170 7194 14172
rect 7218 14170 7274 14172
rect 7298 14170 7354 14172
rect 7058 14118 7104 14170
rect 7104 14118 7114 14170
rect 7138 14118 7168 14170
rect 7168 14118 7180 14170
rect 7180 14118 7194 14170
rect 7218 14118 7232 14170
rect 7232 14118 7244 14170
rect 7244 14118 7274 14170
rect 7298 14118 7308 14170
rect 7308 14118 7354 14170
rect 7058 14116 7114 14118
rect 7138 14116 7194 14118
rect 7218 14116 7274 14118
rect 7298 14116 7354 14118
rect 7058 13082 7114 13084
rect 7138 13082 7194 13084
rect 7218 13082 7274 13084
rect 7298 13082 7354 13084
rect 7058 13030 7104 13082
rect 7104 13030 7114 13082
rect 7138 13030 7168 13082
rect 7168 13030 7180 13082
rect 7180 13030 7194 13082
rect 7218 13030 7232 13082
rect 7232 13030 7244 13082
rect 7244 13030 7274 13082
rect 7298 13030 7308 13082
rect 7308 13030 7354 13082
rect 7058 13028 7114 13030
rect 7138 13028 7194 13030
rect 7218 13028 7274 13030
rect 7298 13028 7354 13030
rect 7058 11994 7114 11996
rect 7138 11994 7194 11996
rect 7218 11994 7274 11996
rect 7298 11994 7354 11996
rect 7058 11942 7104 11994
rect 7104 11942 7114 11994
rect 7138 11942 7168 11994
rect 7168 11942 7180 11994
rect 7180 11942 7194 11994
rect 7218 11942 7232 11994
rect 7232 11942 7244 11994
rect 7244 11942 7274 11994
rect 7298 11942 7308 11994
rect 7308 11942 7354 11994
rect 7058 11940 7114 11942
rect 7138 11940 7194 11942
rect 7218 11940 7274 11942
rect 7298 11940 7354 11942
rect 7058 10906 7114 10908
rect 7138 10906 7194 10908
rect 7218 10906 7274 10908
rect 7298 10906 7354 10908
rect 7058 10854 7104 10906
rect 7104 10854 7114 10906
rect 7138 10854 7168 10906
rect 7168 10854 7180 10906
rect 7180 10854 7194 10906
rect 7218 10854 7232 10906
rect 7232 10854 7244 10906
rect 7244 10854 7274 10906
rect 7298 10854 7308 10906
rect 7308 10854 7354 10906
rect 7058 10852 7114 10854
rect 7138 10852 7194 10854
rect 7218 10852 7274 10854
rect 7298 10852 7354 10854
rect 7058 9818 7114 9820
rect 7138 9818 7194 9820
rect 7218 9818 7274 9820
rect 7298 9818 7354 9820
rect 7058 9766 7104 9818
rect 7104 9766 7114 9818
rect 7138 9766 7168 9818
rect 7168 9766 7180 9818
rect 7180 9766 7194 9818
rect 7218 9766 7232 9818
rect 7232 9766 7244 9818
rect 7244 9766 7274 9818
rect 7298 9766 7308 9818
rect 7308 9766 7354 9818
rect 7058 9764 7114 9766
rect 7138 9764 7194 9766
rect 7218 9764 7274 9766
rect 7298 9764 7354 9766
rect 7058 8730 7114 8732
rect 7138 8730 7194 8732
rect 7218 8730 7274 8732
rect 7298 8730 7354 8732
rect 7058 8678 7104 8730
rect 7104 8678 7114 8730
rect 7138 8678 7168 8730
rect 7168 8678 7180 8730
rect 7180 8678 7194 8730
rect 7218 8678 7232 8730
rect 7232 8678 7244 8730
rect 7244 8678 7274 8730
rect 7298 8678 7308 8730
rect 7308 8678 7354 8730
rect 7058 8676 7114 8678
rect 7138 8676 7194 8678
rect 7218 8676 7274 8678
rect 7298 8676 7354 8678
rect 7058 7642 7114 7644
rect 7138 7642 7194 7644
rect 7218 7642 7274 7644
rect 7298 7642 7354 7644
rect 7058 7590 7104 7642
rect 7104 7590 7114 7642
rect 7138 7590 7168 7642
rect 7168 7590 7180 7642
rect 7180 7590 7194 7642
rect 7218 7590 7232 7642
rect 7232 7590 7244 7642
rect 7244 7590 7274 7642
rect 7298 7590 7308 7642
rect 7308 7590 7354 7642
rect 7058 7588 7114 7590
rect 7138 7588 7194 7590
rect 7218 7588 7274 7590
rect 7298 7588 7354 7590
rect 7058 6554 7114 6556
rect 7138 6554 7194 6556
rect 7218 6554 7274 6556
rect 7298 6554 7354 6556
rect 7058 6502 7104 6554
rect 7104 6502 7114 6554
rect 7138 6502 7168 6554
rect 7168 6502 7180 6554
rect 7180 6502 7194 6554
rect 7218 6502 7232 6554
rect 7232 6502 7244 6554
rect 7244 6502 7274 6554
rect 7298 6502 7308 6554
rect 7308 6502 7354 6554
rect 7058 6500 7114 6502
rect 7138 6500 7194 6502
rect 7218 6500 7274 6502
rect 7298 6500 7354 6502
rect 4007 4922 4063 4924
rect 4087 4922 4143 4924
rect 4167 4922 4223 4924
rect 4247 4922 4303 4924
rect 4007 4870 4053 4922
rect 4053 4870 4063 4922
rect 4087 4870 4117 4922
rect 4117 4870 4129 4922
rect 4129 4870 4143 4922
rect 4167 4870 4181 4922
rect 4181 4870 4193 4922
rect 4193 4870 4223 4922
rect 4247 4870 4257 4922
rect 4257 4870 4303 4922
rect 4007 4868 4063 4870
rect 4087 4868 4143 4870
rect 4167 4868 4223 4870
rect 4247 4868 4303 4870
rect 7058 5466 7114 5468
rect 7138 5466 7194 5468
rect 7218 5466 7274 5468
rect 7298 5466 7354 5468
rect 7058 5414 7104 5466
rect 7104 5414 7114 5466
rect 7138 5414 7168 5466
rect 7168 5414 7180 5466
rect 7180 5414 7194 5466
rect 7218 5414 7232 5466
rect 7232 5414 7244 5466
rect 7244 5414 7274 5466
rect 7298 5414 7308 5466
rect 7308 5414 7354 5466
rect 7058 5412 7114 5414
rect 7138 5412 7194 5414
rect 7218 5412 7274 5414
rect 7298 5412 7354 5414
rect 4007 3834 4063 3836
rect 4087 3834 4143 3836
rect 4167 3834 4223 3836
rect 4247 3834 4303 3836
rect 4007 3782 4053 3834
rect 4053 3782 4063 3834
rect 4087 3782 4117 3834
rect 4117 3782 4129 3834
rect 4129 3782 4143 3834
rect 4167 3782 4181 3834
rect 4181 3782 4193 3834
rect 4193 3782 4223 3834
rect 4247 3782 4257 3834
rect 4257 3782 4303 3834
rect 4007 3780 4063 3782
rect 4087 3780 4143 3782
rect 4167 3780 4223 3782
rect 4247 3780 4303 3782
rect 10110 20154 10166 20156
rect 10190 20154 10246 20156
rect 10270 20154 10326 20156
rect 10350 20154 10406 20156
rect 10110 20102 10156 20154
rect 10156 20102 10166 20154
rect 10190 20102 10220 20154
rect 10220 20102 10232 20154
rect 10232 20102 10246 20154
rect 10270 20102 10284 20154
rect 10284 20102 10296 20154
rect 10296 20102 10326 20154
rect 10350 20102 10360 20154
rect 10360 20102 10406 20154
rect 10110 20100 10166 20102
rect 10190 20100 10246 20102
rect 10270 20100 10326 20102
rect 10350 20100 10406 20102
rect 10110 19066 10166 19068
rect 10190 19066 10246 19068
rect 10270 19066 10326 19068
rect 10350 19066 10406 19068
rect 10110 19014 10156 19066
rect 10156 19014 10166 19066
rect 10190 19014 10220 19066
rect 10220 19014 10232 19066
rect 10232 19014 10246 19066
rect 10270 19014 10284 19066
rect 10284 19014 10296 19066
rect 10296 19014 10326 19066
rect 10350 19014 10360 19066
rect 10360 19014 10406 19066
rect 10110 19012 10166 19014
rect 10190 19012 10246 19014
rect 10270 19012 10326 19014
rect 10350 19012 10406 19014
rect 10110 17978 10166 17980
rect 10190 17978 10246 17980
rect 10270 17978 10326 17980
rect 10350 17978 10406 17980
rect 10110 17926 10156 17978
rect 10156 17926 10166 17978
rect 10190 17926 10220 17978
rect 10220 17926 10232 17978
rect 10232 17926 10246 17978
rect 10270 17926 10284 17978
rect 10284 17926 10296 17978
rect 10296 17926 10326 17978
rect 10350 17926 10360 17978
rect 10360 17926 10406 17978
rect 10110 17924 10166 17926
rect 10190 17924 10246 17926
rect 10270 17924 10326 17926
rect 10350 17924 10406 17926
rect 10110 16890 10166 16892
rect 10190 16890 10246 16892
rect 10270 16890 10326 16892
rect 10350 16890 10406 16892
rect 10110 16838 10156 16890
rect 10156 16838 10166 16890
rect 10190 16838 10220 16890
rect 10220 16838 10232 16890
rect 10232 16838 10246 16890
rect 10270 16838 10284 16890
rect 10284 16838 10296 16890
rect 10296 16838 10326 16890
rect 10350 16838 10360 16890
rect 10360 16838 10406 16890
rect 10110 16836 10166 16838
rect 10190 16836 10246 16838
rect 10270 16836 10326 16838
rect 10350 16836 10406 16838
rect 10110 15802 10166 15804
rect 10190 15802 10246 15804
rect 10270 15802 10326 15804
rect 10350 15802 10406 15804
rect 10110 15750 10156 15802
rect 10156 15750 10166 15802
rect 10190 15750 10220 15802
rect 10220 15750 10232 15802
rect 10232 15750 10246 15802
rect 10270 15750 10284 15802
rect 10284 15750 10296 15802
rect 10296 15750 10326 15802
rect 10350 15750 10360 15802
rect 10360 15750 10406 15802
rect 10110 15748 10166 15750
rect 10190 15748 10246 15750
rect 10270 15748 10326 15750
rect 10350 15748 10406 15750
rect 10110 14714 10166 14716
rect 10190 14714 10246 14716
rect 10270 14714 10326 14716
rect 10350 14714 10406 14716
rect 10110 14662 10156 14714
rect 10156 14662 10166 14714
rect 10190 14662 10220 14714
rect 10220 14662 10232 14714
rect 10232 14662 10246 14714
rect 10270 14662 10284 14714
rect 10284 14662 10296 14714
rect 10296 14662 10326 14714
rect 10350 14662 10360 14714
rect 10360 14662 10406 14714
rect 10110 14660 10166 14662
rect 10190 14660 10246 14662
rect 10270 14660 10326 14662
rect 10350 14660 10406 14662
rect 10110 13626 10166 13628
rect 10190 13626 10246 13628
rect 10270 13626 10326 13628
rect 10350 13626 10406 13628
rect 10110 13574 10156 13626
rect 10156 13574 10166 13626
rect 10190 13574 10220 13626
rect 10220 13574 10232 13626
rect 10232 13574 10246 13626
rect 10270 13574 10284 13626
rect 10284 13574 10296 13626
rect 10296 13574 10326 13626
rect 10350 13574 10360 13626
rect 10360 13574 10406 13626
rect 10110 13572 10166 13574
rect 10190 13572 10246 13574
rect 10270 13572 10326 13574
rect 10350 13572 10406 13574
rect 10110 12538 10166 12540
rect 10190 12538 10246 12540
rect 10270 12538 10326 12540
rect 10350 12538 10406 12540
rect 10110 12486 10156 12538
rect 10156 12486 10166 12538
rect 10190 12486 10220 12538
rect 10220 12486 10232 12538
rect 10232 12486 10246 12538
rect 10270 12486 10284 12538
rect 10284 12486 10296 12538
rect 10296 12486 10326 12538
rect 10350 12486 10360 12538
rect 10360 12486 10406 12538
rect 10110 12484 10166 12486
rect 10190 12484 10246 12486
rect 10270 12484 10326 12486
rect 10350 12484 10406 12486
rect 10110 11450 10166 11452
rect 10190 11450 10246 11452
rect 10270 11450 10326 11452
rect 10350 11450 10406 11452
rect 10110 11398 10156 11450
rect 10156 11398 10166 11450
rect 10190 11398 10220 11450
rect 10220 11398 10232 11450
rect 10232 11398 10246 11450
rect 10270 11398 10284 11450
rect 10284 11398 10296 11450
rect 10296 11398 10326 11450
rect 10350 11398 10360 11450
rect 10360 11398 10406 11450
rect 10110 11396 10166 11398
rect 10190 11396 10246 11398
rect 10270 11396 10326 11398
rect 10350 11396 10406 11398
rect 13161 19610 13217 19612
rect 13241 19610 13297 19612
rect 13321 19610 13377 19612
rect 13401 19610 13457 19612
rect 13161 19558 13207 19610
rect 13207 19558 13217 19610
rect 13241 19558 13271 19610
rect 13271 19558 13283 19610
rect 13283 19558 13297 19610
rect 13321 19558 13335 19610
rect 13335 19558 13347 19610
rect 13347 19558 13377 19610
rect 13401 19558 13411 19610
rect 13411 19558 13457 19610
rect 13161 19556 13217 19558
rect 13241 19556 13297 19558
rect 13321 19556 13377 19558
rect 13401 19556 13457 19558
rect 13161 18522 13217 18524
rect 13241 18522 13297 18524
rect 13321 18522 13377 18524
rect 13401 18522 13457 18524
rect 13161 18470 13207 18522
rect 13207 18470 13217 18522
rect 13241 18470 13271 18522
rect 13271 18470 13283 18522
rect 13283 18470 13297 18522
rect 13321 18470 13335 18522
rect 13335 18470 13347 18522
rect 13347 18470 13377 18522
rect 13401 18470 13411 18522
rect 13411 18470 13457 18522
rect 13161 18468 13217 18470
rect 13241 18468 13297 18470
rect 13321 18468 13377 18470
rect 13401 18468 13457 18470
rect 13161 17434 13217 17436
rect 13241 17434 13297 17436
rect 13321 17434 13377 17436
rect 13401 17434 13457 17436
rect 13161 17382 13207 17434
rect 13207 17382 13217 17434
rect 13241 17382 13271 17434
rect 13271 17382 13283 17434
rect 13283 17382 13297 17434
rect 13321 17382 13335 17434
rect 13335 17382 13347 17434
rect 13347 17382 13377 17434
rect 13401 17382 13411 17434
rect 13411 17382 13457 17434
rect 13161 17380 13217 17382
rect 13241 17380 13297 17382
rect 13321 17380 13377 17382
rect 13401 17380 13457 17382
rect 13161 16346 13217 16348
rect 13241 16346 13297 16348
rect 13321 16346 13377 16348
rect 13401 16346 13457 16348
rect 13161 16294 13207 16346
rect 13207 16294 13217 16346
rect 13241 16294 13271 16346
rect 13271 16294 13283 16346
rect 13283 16294 13297 16346
rect 13321 16294 13335 16346
rect 13335 16294 13347 16346
rect 13347 16294 13377 16346
rect 13401 16294 13411 16346
rect 13411 16294 13457 16346
rect 13161 16292 13217 16294
rect 13241 16292 13297 16294
rect 13321 16292 13377 16294
rect 13401 16292 13457 16294
rect 13161 15258 13217 15260
rect 13241 15258 13297 15260
rect 13321 15258 13377 15260
rect 13401 15258 13457 15260
rect 13161 15206 13207 15258
rect 13207 15206 13217 15258
rect 13241 15206 13271 15258
rect 13271 15206 13283 15258
rect 13283 15206 13297 15258
rect 13321 15206 13335 15258
rect 13335 15206 13347 15258
rect 13347 15206 13377 15258
rect 13401 15206 13411 15258
rect 13411 15206 13457 15258
rect 13161 15204 13217 15206
rect 13241 15204 13297 15206
rect 13321 15204 13377 15206
rect 13401 15204 13457 15206
rect 13161 14170 13217 14172
rect 13241 14170 13297 14172
rect 13321 14170 13377 14172
rect 13401 14170 13457 14172
rect 13161 14118 13207 14170
rect 13207 14118 13217 14170
rect 13241 14118 13271 14170
rect 13271 14118 13283 14170
rect 13283 14118 13297 14170
rect 13321 14118 13335 14170
rect 13335 14118 13347 14170
rect 13347 14118 13377 14170
rect 13401 14118 13411 14170
rect 13411 14118 13457 14170
rect 13161 14116 13217 14118
rect 13241 14116 13297 14118
rect 13321 14116 13377 14118
rect 13401 14116 13457 14118
rect 13161 13082 13217 13084
rect 13241 13082 13297 13084
rect 13321 13082 13377 13084
rect 13401 13082 13457 13084
rect 13161 13030 13207 13082
rect 13207 13030 13217 13082
rect 13241 13030 13271 13082
rect 13271 13030 13283 13082
rect 13283 13030 13297 13082
rect 13321 13030 13335 13082
rect 13335 13030 13347 13082
rect 13347 13030 13377 13082
rect 13401 13030 13411 13082
rect 13411 13030 13457 13082
rect 13161 13028 13217 13030
rect 13241 13028 13297 13030
rect 13321 13028 13377 13030
rect 13401 13028 13457 13030
rect 13161 11994 13217 11996
rect 13241 11994 13297 11996
rect 13321 11994 13377 11996
rect 13401 11994 13457 11996
rect 13161 11942 13207 11994
rect 13207 11942 13217 11994
rect 13241 11942 13271 11994
rect 13271 11942 13283 11994
rect 13283 11942 13297 11994
rect 13321 11942 13335 11994
rect 13335 11942 13347 11994
rect 13347 11942 13377 11994
rect 13401 11942 13411 11994
rect 13411 11942 13457 11994
rect 13161 11940 13217 11942
rect 13241 11940 13297 11942
rect 13321 11940 13377 11942
rect 13401 11940 13457 11942
rect 10110 10362 10166 10364
rect 10190 10362 10246 10364
rect 10270 10362 10326 10364
rect 10350 10362 10406 10364
rect 10110 10310 10156 10362
rect 10156 10310 10166 10362
rect 10190 10310 10220 10362
rect 10220 10310 10232 10362
rect 10232 10310 10246 10362
rect 10270 10310 10284 10362
rect 10284 10310 10296 10362
rect 10296 10310 10326 10362
rect 10350 10310 10360 10362
rect 10360 10310 10406 10362
rect 10110 10308 10166 10310
rect 10190 10308 10246 10310
rect 10270 10308 10326 10310
rect 10350 10308 10406 10310
rect 10110 9274 10166 9276
rect 10190 9274 10246 9276
rect 10270 9274 10326 9276
rect 10350 9274 10406 9276
rect 10110 9222 10156 9274
rect 10156 9222 10166 9274
rect 10190 9222 10220 9274
rect 10220 9222 10232 9274
rect 10232 9222 10246 9274
rect 10270 9222 10284 9274
rect 10284 9222 10296 9274
rect 10296 9222 10326 9274
rect 10350 9222 10360 9274
rect 10360 9222 10406 9274
rect 10110 9220 10166 9222
rect 10190 9220 10246 9222
rect 10270 9220 10326 9222
rect 10350 9220 10406 9222
rect 10110 8186 10166 8188
rect 10190 8186 10246 8188
rect 10270 8186 10326 8188
rect 10350 8186 10406 8188
rect 10110 8134 10156 8186
rect 10156 8134 10166 8186
rect 10190 8134 10220 8186
rect 10220 8134 10232 8186
rect 10232 8134 10246 8186
rect 10270 8134 10284 8186
rect 10284 8134 10296 8186
rect 10296 8134 10326 8186
rect 10350 8134 10360 8186
rect 10360 8134 10406 8186
rect 10110 8132 10166 8134
rect 10190 8132 10246 8134
rect 10270 8132 10326 8134
rect 10350 8132 10406 8134
rect 7058 4378 7114 4380
rect 7138 4378 7194 4380
rect 7218 4378 7274 4380
rect 7298 4378 7354 4380
rect 7058 4326 7104 4378
rect 7104 4326 7114 4378
rect 7138 4326 7168 4378
rect 7168 4326 7180 4378
rect 7180 4326 7194 4378
rect 7218 4326 7232 4378
rect 7232 4326 7244 4378
rect 7244 4326 7274 4378
rect 7298 4326 7308 4378
rect 7308 4326 7354 4378
rect 7058 4324 7114 4326
rect 7138 4324 7194 4326
rect 7218 4324 7274 4326
rect 7298 4324 7354 4326
rect 10110 7098 10166 7100
rect 10190 7098 10246 7100
rect 10270 7098 10326 7100
rect 10350 7098 10406 7100
rect 10110 7046 10156 7098
rect 10156 7046 10166 7098
rect 10190 7046 10220 7098
rect 10220 7046 10232 7098
rect 10232 7046 10246 7098
rect 10270 7046 10284 7098
rect 10284 7046 10296 7098
rect 10296 7046 10326 7098
rect 10350 7046 10360 7098
rect 10360 7046 10406 7098
rect 10110 7044 10166 7046
rect 10190 7044 10246 7046
rect 10270 7044 10326 7046
rect 10350 7044 10406 7046
rect 10110 6010 10166 6012
rect 10190 6010 10246 6012
rect 10270 6010 10326 6012
rect 10350 6010 10406 6012
rect 10110 5958 10156 6010
rect 10156 5958 10166 6010
rect 10190 5958 10220 6010
rect 10220 5958 10232 6010
rect 10232 5958 10246 6010
rect 10270 5958 10284 6010
rect 10284 5958 10296 6010
rect 10296 5958 10326 6010
rect 10350 5958 10360 6010
rect 10360 5958 10406 6010
rect 10110 5956 10166 5958
rect 10190 5956 10246 5958
rect 10270 5956 10326 5958
rect 10350 5956 10406 5958
rect 7058 3290 7114 3292
rect 7138 3290 7194 3292
rect 7218 3290 7274 3292
rect 7298 3290 7354 3292
rect 7058 3238 7104 3290
rect 7104 3238 7114 3290
rect 7138 3238 7168 3290
rect 7168 3238 7180 3290
rect 7180 3238 7194 3290
rect 7218 3238 7232 3290
rect 7232 3238 7244 3290
rect 7244 3238 7274 3290
rect 7298 3238 7308 3290
rect 7308 3238 7354 3290
rect 7058 3236 7114 3238
rect 7138 3236 7194 3238
rect 7218 3236 7274 3238
rect 7298 3236 7354 3238
rect 10110 4922 10166 4924
rect 10190 4922 10246 4924
rect 10270 4922 10326 4924
rect 10350 4922 10406 4924
rect 10110 4870 10156 4922
rect 10156 4870 10166 4922
rect 10190 4870 10220 4922
rect 10220 4870 10232 4922
rect 10232 4870 10246 4922
rect 10270 4870 10284 4922
rect 10284 4870 10296 4922
rect 10296 4870 10326 4922
rect 10350 4870 10360 4922
rect 10360 4870 10406 4922
rect 10110 4868 10166 4870
rect 10190 4868 10246 4870
rect 10270 4868 10326 4870
rect 10350 4868 10406 4870
rect 10110 3834 10166 3836
rect 10190 3834 10246 3836
rect 10270 3834 10326 3836
rect 10350 3834 10406 3836
rect 10110 3782 10156 3834
rect 10156 3782 10166 3834
rect 10190 3782 10220 3834
rect 10220 3782 10232 3834
rect 10232 3782 10246 3834
rect 10270 3782 10284 3834
rect 10284 3782 10296 3834
rect 10296 3782 10326 3834
rect 10350 3782 10360 3834
rect 10360 3782 10406 3834
rect 10110 3780 10166 3782
rect 10190 3780 10246 3782
rect 10270 3780 10326 3782
rect 10350 3780 10406 3782
rect 13161 10906 13217 10908
rect 13241 10906 13297 10908
rect 13321 10906 13377 10908
rect 13401 10906 13457 10908
rect 13161 10854 13207 10906
rect 13207 10854 13217 10906
rect 13241 10854 13271 10906
rect 13271 10854 13283 10906
rect 13283 10854 13297 10906
rect 13321 10854 13335 10906
rect 13335 10854 13347 10906
rect 13347 10854 13377 10906
rect 13401 10854 13411 10906
rect 13411 10854 13457 10906
rect 13161 10852 13217 10854
rect 13241 10852 13297 10854
rect 13321 10852 13377 10854
rect 13401 10852 13457 10854
rect 13161 9818 13217 9820
rect 13241 9818 13297 9820
rect 13321 9818 13377 9820
rect 13401 9818 13457 9820
rect 13161 9766 13207 9818
rect 13207 9766 13217 9818
rect 13241 9766 13271 9818
rect 13271 9766 13283 9818
rect 13283 9766 13297 9818
rect 13321 9766 13335 9818
rect 13335 9766 13347 9818
rect 13347 9766 13377 9818
rect 13401 9766 13411 9818
rect 13411 9766 13457 9818
rect 13161 9764 13217 9766
rect 13241 9764 13297 9766
rect 13321 9764 13377 9766
rect 13401 9764 13457 9766
rect 13161 8730 13217 8732
rect 13241 8730 13297 8732
rect 13321 8730 13377 8732
rect 13401 8730 13457 8732
rect 13161 8678 13207 8730
rect 13207 8678 13217 8730
rect 13241 8678 13271 8730
rect 13271 8678 13283 8730
rect 13283 8678 13297 8730
rect 13321 8678 13335 8730
rect 13335 8678 13347 8730
rect 13347 8678 13377 8730
rect 13401 8678 13411 8730
rect 13411 8678 13457 8730
rect 13161 8676 13217 8678
rect 13241 8676 13297 8678
rect 13321 8676 13377 8678
rect 13401 8676 13457 8678
rect 13161 7642 13217 7644
rect 13241 7642 13297 7644
rect 13321 7642 13377 7644
rect 13401 7642 13457 7644
rect 13161 7590 13207 7642
rect 13207 7590 13217 7642
rect 13241 7590 13271 7642
rect 13271 7590 13283 7642
rect 13283 7590 13297 7642
rect 13321 7590 13335 7642
rect 13335 7590 13347 7642
rect 13347 7590 13377 7642
rect 13401 7590 13411 7642
rect 13411 7590 13457 7642
rect 13161 7588 13217 7590
rect 13241 7588 13297 7590
rect 13321 7588 13377 7590
rect 13401 7588 13457 7590
rect 13161 6554 13217 6556
rect 13241 6554 13297 6556
rect 13321 6554 13377 6556
rect 13401 6554 13457 6556
rect 13161 6502 13207 6554
rect 13207 6502 13217 6554
rect 13241 6502 13271 6554
rect 13271 6502 13283 6554
rect 13283 6502 13297 6554
rect 13321 6502 13335 6554
rect 13335 6502 13347 6554
rect 13347 6502 13377 6554
rect 13401 6502 13411 6554
rect 13411 6502 13457 6554
rect 13161 6500 13217 6502
rect 13241 6500 13297 6502
rect 13321 6500 13377 6502
rect 13401 6500 13457 6502
rect 13161 5466 13217 5468
rect 13241 5466 13297 5468
rect 13321 5466 13377 5468
rect 13401 5466 13457 5468
rect 13161 5414 13207 5466
rect 13207 5414 13217 5466
rect 13241 5414 13271 5466
rect 13271 5414 13283 5466
rect 13283 5414 13297 5466
rect 13321 5414 13335 5466
rect 13335 5414 13347 5466
rect 13347 5414 13377 5466
rect 13401 5414 13411 5466
rect 13411 5414 13457 5466
rect 13161 5412 13217 5414
rect 13241 5412 13297 5414
rect 13321 5412 13377 5414
rect 13401 5412 13457 5414
rect 16212 20154 16268 20156
rect 16292 20154 16348 20156
rect 16372 20154 16428 20156
rect 16452 20154 16508 20156
rect 16212 20102 16258 20154
rect 16258 20102 16268 20154
rect 16292 20102 16322 20154
rect 16322 20102 16334 20154
rect 16334 20102 16348 20154
rect 16372 20102 16386 20154
rect 16386 20102 16398 20154
rect 16398 20102 16428 20154
rect 16452 20102 16462 20154
rect 16462 20102 16508 20154
rect 16212 20100 16268 20102
rect 16292 20100 16348 20102
rect 16372 20100 16428 20102
rect 16452 20100 16508 20102
rect 16212 19066 16268 19068
rect 16292 19066 16348 19068
rect 16372 19066 16428 19068
rect 16452 19066 16508 19068
rect 16212 19014 16258 19066
rect 16258 19014 16268 19066
rect 16292 19014 16322 19066
rect 16322 19014 16334 19066
rect 16334 19014 16348 19066
rect 16372 19014 16386 19066
rect 16386 19014 16398 19066
rect 16398 19014 16428 19066
rect 16452 19014 16462 19066
rect 16462 19014 16508 19066
rect 16212 19012 16268 19014
rect 16292 19012 16348 19014
rect 16372 19012 16428 19014
rect 16452 19012 16508 19014
rect 16212 17978 16268 17980
rect 16292 17978 16348 17980
rect 16372 17978 16428 17980
rect 16452 17978 16508 17980
rect 16212 17926 16258 17978
rect 16258 17926 16268 17978
rect 16292 17926 16322 17978
rect 16322 17926 16334 17978
rect 16334 17926 16348 17978
rect 16372 17926 16386 17978
rect 16386 17926 16398 17978
rect 16398 17926 16428 17978
rect 16452 17926 16462 17978
rect 16462 17926 16508 17978
rect 16212 17924 16268 17926
rect 16292 17924 16348 17926
rect 16372 17924 16428 17926
rect 16452 17924 16508 17926
rect 16212 16890 16268 16892
rect 16292 16890 16348 16892
rect 16372 16890 16428 16892
rect 16452 16890 16508 16892
rect 16212 16838 16258 16890
rect 16258 16838 16268 16890
rect 16292 16838 16322 16890
rect 16322 16838 16334 16890
rect 16334 16838 16348 16890
rect 16372 16838 16386 16890
rect 16386 16838 16398 16890
rect 16398 16838 16428 16890
rect 16452 16838 16462 16890
rect 16462 16838 16508 16890
rect 16212 16836 16268 16838
rect 16292 16836 16348 16838
rect 16372 16836 16428 16838
rect 16452 16836 16508 16838
rect 16212 15802 16268 15804
rect 16292 15802 16348 15804
rect 16372 15802 16428 15804
rect 16452 15802 16508 15804
rect 16212 15750 16258 15802
rect 16258 15750 16268 15802
rect 16292 15750 16322 15802
rect 16322 15750 16334 15802
rect 16334 15750 16348 15802
rect 16372 15750 16386 15802
rect 16386 15750 16398 15802
rect 16398 15750 16428 15802
rect 16452 15750 16462 15802
rect 16462 15750 16508 15802
rect 16212 15748 16268 15750
rect 16292 15748 16348 15750
rect 16372 15748 16428 15750
rect 16452 15748 16508 15750
rect 16212 14714 16268 14716
rect 16292 14714 16348 14716
rect 16372 14714 16428 14716
rect 16452 14714 16508 14716
rect 16212 14662 16258 14714
rect 16258 14662 16268 14714
rect 16292 14662 16322 14714
rect 16322 14662 16334 14714
rect 16334 14662 16348 14714
rect 16372 14662 16386 14714
rect 16386 14662 16398 14714
rect 16398 14662 16428 14714
rect 16452 14662 16462 14714
rect 16462 14662 16508 14714
rect 16212 14660 16268 14662
rect 16292 14660 16348 14662
rect 16372 14660 16428 14662
rect 16452 14660 16508 14662
rect 16212 13626 16268 13628
rect 16292 13626 16348 13628
rect 16372 13626 16428 13628
rect 16452 13626 16508 13628
rect 16212 13574 16258 13626
rect 16258 13574 16268 13626
rect 16292 13574 16322 13626
rect 16322 13574 16334 13626
rect 16334 13574 16348 13626
rect 16372 13574 16386 13626
rect 16386 13574 16398 13626
rect 16398 13574 16428 13626
rect 16452 13574 16462 13626
rect 16462 13574 16508 13626
rect 16212 13572 16268 13574
rect 16292 13572 16348 13574
rect 16372 13572 16428 13574
rect 16452 13572 16508 13574
rect 16212 12538 16268 12540
rect 16292 12538 16348 12540
rect 16372 12538 16428 12540
rect 16452 12538 16508 12540
rect 16212 12486 16258 12538
rect 16258 12486 16268 12538
rect 16292 12486 16322 12538
rect 16322 12486 16334 12538
rect 16334 12486 16348 12538
rect 16372 12486 16386 12538
rect 16386 12486 16398 12538
rect 16398 12486 16428 12538
rect 16452 12486 16462 12538
rect 16462 12486 16508 12538
rect 16212 12484 16268 12486
rect 16292 12484 16348 12486
rect 16372 12484 16428 12486
rect 16452 12484 16508 12486
rect 15842 11192 15898 11248
rect 16212 11450 16268 11452
rect 16292 11450 16348 11452
rect 16372 11450 16428 11452
rect 16452 11450 16508 11452
rect 16212 11398 16258 11450
rect 16258 11398 16268 11450
rect 16292 11398 16322 11450
rect 16322 11398 16334 11450
rect 16334 11398 16348 11450
rect 16372 11398 16386 11450
rect 16386 11398 16398 11450
rect 16398 11398 16428 11450
rect 16452 11398 16462 11450
rect 16462 11398 16508 11450
rect 16212 11396 16268 11398
rect 16292 11396 16348 11398
rect 16372 11396 16428 11398
rect 16452 11396 16508 11398
rect 16212 10362 16268 10364
rect 16292 10362 16348 10364
rect 16372 10362 16428 10364
rect 16452 10362 16508 10364
rect 16212 10310 16258 10362
rect 16258 10310 16268 10362
rect 16292 10310 16322 10362
rect 16322 10310 16334 10362
rect 16334 10310 16348 10362
rect 16372 10310 16386 10362
rect 16386 10310 16398 10362
rect 16398 10310 16428 10362
rect 16452 10310 16462 10362
rect 16462 10310 16508 10362
rect 16212 10308 16268 10310
rect 16292 10308 16348 10310
rect 16372 10308 16428 10310
rect 16452 10308 16508 10310
rect 16212 9274 16268 9276
rect 16292 9274 16348 9276
rect 16372 9274 16428 9276
rect 16452 9274 16508 9276
rect 16212 9222 16258 9274
rect 16258 9222 16268 9274
rect 16292 9222 16322 9274
rect 16322 9222 16334 9274
rect 16334 9222 16348 9274
rect 16372 9222 16386 9274
rect 16386 9222 16398 9274
rect 16398 9222 16428 9274
rect 16452 9222 16462 9274
rect 16462 9222 16508 9274
rect 16212 9220 16268 9222
rect 16292 9220 16348 9222
rect 16372 9220 16428 9222
rect 16452 9220 16508 9222
rect 16212 8186 16268 8188
rect 16292 8186 16348 8188
rect 16372 8186 16428 8188
rect 16452 8186 16508 8188
rect 16212 8134 16258 8186
rect 16258 8134 16268 8186
rect 16292 8134 16322 8186
rect 16322 8134 16334 8186
rect 16334 8134 16348 8186
rect 16372 8134 16386 8186
rect 16386 8134 16398 8186
rect 16398 8134 16428 8186
rect 16452 8134 16462 8186
rect 16462 8134 16508 8186
rect 16212 8132 16268 8134
rect 16292 8132 16348 8134
rect 16372 8132 16428 8134
rect 16452 8132 16508 8134
rect 16212 7098 16268 7100
rect 16292 7098 16348 7100
rect 16372 7098 16428 7100
rect 16452 7098 16508 7100
rect 16212 7046 16258 7098
rect 16258 7046 16268 7098
rect 16292 7046 16322 7098
rect 16322 7046 16334 7098
rect 16334 7046 16348 7098
rect 16372 7046 16386 7098
rect 16386 7046 16398 7098
rect 16398 7046 16428 7098
rect 16452 7046 16462 7098
rect 16462 7046 16508 7098
rect 16212 7044 16268 7046
rect 16292 7044 16348 7046
rect 16372 7044 16428 7046
rect 16452 7044 16508 7046
rect 13161 4378 13217 4380
rect 13241 4378 13297 4380
rect 13321 4378 13377 4380
rect 13401 4378 13457 4380
rect 13161 4326 13207 4378
rect 13207 4326 13217 4378
rect 13241 4326 13271 4378
rect 13271 4326 13283 4378
rect 13283 4326 13297 4378
rect 13321 4326 13335 4378
rect 13335 4326 13347 4378
rect 13347 4326 13377 4378
rect 13401 4326 13411 4378
rect 13411 4326 13457 4378
rect 13161 4324 13217 4326
rect 13241 4324 13297 4326
rect 13321 4324 13377 4326
rect 13401 4324 13457 4326
rect 13161 3290 13217 3292
rect 13241 3290 13297 3292
rect 13321 3290 13377 3292
rect 13401 3290 13457 3292
rect 13161 3238 13207 3290
rect 13207 3238 13217 3290
rect 13241 3238 13271 3290
rect 13271 3238 13283 3290
rect 13283 3238 13297 3290
rect 13321 3238 13335 3290
rect 13335 3238 13347 3290
rect 13347 3238 13377 3290
rect 13401 3238 13411 3290
rect 13411 3238 13457 3290
rect 13161 3236 13217 3238
rect 13241 3236 13297 3238
rect 13321 3236 13377 3238
rect 13401 3236 13457 3238
rect 16212 6010 16268 6012
rect 16292 6010 16348 6012
rect 16372 6010 16428 6012
rect 16452 6010 16508 6012
rect 16212 5958 16258 6010
rect 16258 5958 16268 6010
rect 16292 5958 16322 6010
rect 16322 5958 16334 6010
rect 16334 5958 16348 6010
rect 16372 5958 16386 6010
rect 16386 5958 16398 6010
rect 16398 5958 16428 6010
rect 16452 5958 16462 6010
rect 16462 5958 16508 6010
rect 16212 5956 16268 5958
rect 16292 5956 16348 5958
rect 16372 5956 16428 5958
rect 16452 5956 16508 5958
rect 16212 4922 16268 4924
rect 16292 4922 16348 4924
rect 16372 4922 16428 4924
rect 16452 4922 16508 4924
rect 16212 4870 16258 4922
rect 16258 4870 16268 4922
rect 16292 4870 16322 4922
rect 16322 4870 16334 4922
rect 16334 4870 16348 4922
rect 16372 4870 16386 4922
rect 16386 4870 16398 4922
rect 16398 4870 16428 4922
rect 16452 4870 16462 4922
rect 16462 4870 16508 4922
rect 16212 4868 16268 4870
rect 16292 4868 16348 4870
rect 16372 4868 16428 4870
rect 16452 4868 16508 4870
rect 16212 3834 16268 3836
rect 16292 3834 16348 3836
rect 16372 3834 16428 3836
rect 16452 3834 16508 3836
rect 16212 3782 16258 3834
rect 16258 3782 16268 3834
rect 16292 3782 16322 3834
rect 16322 3782 16334 3834
rect 16334 3782 16348 3834
rect 16372 3782 16386 3834
rect 16386 3782 16398 3834
rect 16398 3782 16428 3834
rect 16452 3782 16462 3834
rect 16462 3782 16508 3834
rect 16212 3780 16268 3782
rect 16292 3780 16348 3782
rect 16372 3780 16428 3782
rect 16452 3780 16508 3782
rect 4007 2746 4063 2748
rect 4087 2746 4143 2748
rect 4167 2746 4223 2748
rect 4247 2746 4303 2748
rect 4007 2694 4053 2746
rect 4053 2694 4063 2746
rect 4087 2694 4117 2746
rect 4117 2694 4129 2746
rect 4129 2694 4143 2746
rect 4167 2694 4181 2746
rect 4181 2694 4193 2746
rect 4193 2694 4223 2746
rect 4247 2694 4257 2746
rect 4257 2694 4303 2746
rect 4007 2692 4063 2694
rect 4087 2692 4143 2694
rect 4167 2692 4223 2694
rect 4247 2692 4303 2694
rect 10110 2746 10166 2748
rect 10190 2746 10246 2748
rect 10270 2746 10326 2748
rect 10350 2746 10406 2748
rect 10110 2694 10156 2746
rect 10156 2694 10166 2746
rect 10190 2694 10220 2746
rect 10220 2694 10232 2746
rect 10232 2694 10246 2746
rect 10270 2694 10284 2746
rect 10284 2694 10296 2746
rect 10296 2694 10326 2746
rect 10350 2694 10360 2746
rect 10360 2694 10406 2746
rect 10110 2692 10166 2694
rect 10190 2692 10246 2694
rect 10270 2692 10326 2694
rect 10350 2692 10406 2694
rect 16212 2746 16268 2748
rect 16292 2746 16348 2748
rect 16372 2746 16428 2748
rect 16452 2746 16508 2748
rect 16212 2694 16258 2746
rect 16258 2694 16268 2746
rect 16292 2694 16322 2746
rect 16322 2694 16334 2746
rect 16334 2694 16348 2746
rect 16372 2694 16386 2746
rect 16386 2694 16398 2746
rect 16398 2694 16428 2746
rect 16452 2694 16462 2746
rect 16462 2694 16508 2746
rect 16212 2692 16268 2694
rect 16292 2692 16348 2694
rect 16372 2692 16428 2694
rect 16452 2692 16508 2694
rect 7058 2202 7114 2204
rect 7138 2202 7194 2204
rect 7218 2202 7274 2204
rect 7298 2202 7354 2204
rect 7058 2150 7104 2202
rect 7104 2150 7114 2202
rect 7138 2150 7168 2202
rect 7168 2150 7180 2202
rect 7180 2150 7194 2202
rect 7218 2150 7232 2202
rect 7232 2150 7244 2202
rect 7244 2150 7274 2202
rect 7298 2150 7308 2202
rect 7308 2150 7354 2202
rect 7058 2148 7114 2150
rect 7138 2148 7194 2150
rect 7218 2148 7274 2150
rect 7298 2148 7354 2150
rect 13161 2202 13217 2204
rect 13241 2202 13297 2204
rect 13321 2202 13377 2204
rect 13401 2202 13457 2204
rect 13161 2150 13207 2202
rect 13207 2150 13217 2202
rect 13241 2150 13271 2202
rect 13271 2150 13283 2202
rect 13283 2150 13297 2202
rect 13321 2150 13335 2202
rect 13335 2150 13347 2202
rect 13347 2150 13377 2202
rect 13401 2150 13411 2202
rect 13411 2150 13457 2202
rect 13161 2148 13217 2150
rect 13241 2148 13297 2150
rect 13321 2148 13377 2150
rect 13401 2148 13457 2150
<< metal3 >>
rect 3995 20160 4315 20161
rect 3995 20096 4003 20160
rect 4067 20096 4083 20160
rect 4147 20096 4163 20160
rect 4227 20096 4243 20160
rect 4307 20096 4315 20160
rect 3995 20095 4315 20096
rect 10098 20160 10418 20161
rect 10098 20096 10106 20160
rect 10170 20096 10186 20160
rect 10250 20096 10266 20160
rect 10330 20096 10346 20160
rect 10410 20096 10418 20160
rect 10098 20095 10418 20096
rect 16200 20160 16520 20161
rect 16200 20096 16208 20160
rect 16272 20096 16288 20160
rect 16352 20096 16368 20160
rect 16432 20096 16448 20160
rect 16512 20096 16520 20160
rect 16200 20095 16520 20096
rect 7046 19616 7366 19617
rect 7046 19552 7054 19616
rect 7118 19552 7134 19616
rect 7198 19552 7214 19616
rect 7278 19552 7294 19616
rect 7358 19552 7366 19616
rect 7046 19551 7366 19552
rect 13149 19616 13469 19617
rect 13149 19552 13157 19616
rect 13221 19552 13237 19616
rect 13301 19552 13317 19616
rect 13381 19552 13397 19616
rect 13461 19552 13469 19616
rect 13149 19551 13469 19552
rect 3995 19072 4315 19073
rect 3995 19008 4003 19072
rect 4067 19008 4083 19072
rect 4147 19008 4163 19072
rect 4227 19008 4243 19072
rect 4307 19008 4315 19072
rect 3995 19007 4315 19008
rect 10098 19072 10418 19073
rect 10098 19008 10106 19072
rect 10170 19008 10186 19072
rect 10250 19008 10266 19072
rect 10330 19008 10346 19072
rect 10410 19008 10418 19072
rect 10098 19007 10418 19008
rect 16200 19072 16520 19073
rect 16200 19008 16208 19072
rect 16272 19008 16288 19072
rect 16352 19008 16368 19072
rect 16432 19008 16448 19072
rect 16512 19008 16520 19072
rect 16200 19007 16520 19008
rect 7046 18528 7366 18529
rect 7046 18464 7054 18528
rect 7118 18464 7134 18528
rect 7198 18464 7214 18528
rect 7278 18464 7294 18528
rect 7358 18464 7366 18528
rect 7046 18463 7366 18464
rect 13149 18528 13469 18529
rect 13149 18464 13157 18528
rect 13221 18464 13237 18528
rect 13301 18464 13317 18528
rect 13381 18464 13397 18528
rect 13461 18464 13469 18528
rect 13149 18463 13469 18464
rect 3995 17984 4315 17985
rect 3995 17920 4003 17984
rect 4067 17920 4083 17984
rect 4147 17920 4163 17984
rect 4227 17920 4243 17984
rect 4307 17920 4315 17984
rect 3995 17919 4315 17920
rect 10098 17984 10418 17985
rect 10098 17920 10106 17984
rect 10170 17920 10186 17984
rect 10250 17920 10266 17984
rect 10330 17920 10346 17984
rect 10410 17920 10418 17984
rect 10098 17919 10418 17920
rect 16200 17984 16520 17985
rect 16200 17920 16208 17984
rect 16272 17920 16288 17984
rect 16352 17920 16368 17984
rect 16432 17920 16448 17984
rect 16512 17920 16520 17984
rect 16200 17919 16520 17920
rect 7046 17440 7366 17441
rect 7046 17376 7054 17440
rect 7118 17376 7134 17440
rect 7198 17376 7214 17440
rect 7278 17376 7294 17440
rect 7358 17376 7366 17440
rect 7046 17375 7366 17376
rect 13149 17440 13469 17441
rect 13149 17376 13157 17440
rect 13221 17376 13237 17440
rect 13301 17376 13317 17440
rect 13381 17376 13397 17440
rect 13461 17376 13469 17440
rect 13149 17375 13469 17376
rect 3995 16896 4315 16897
rect 3995 16832 4003 16896
rect 4067 16832 4083 16896
rect 4147 16832 4163 16896
rect 4227 16832 4243 16896
rect 4307 16832 4315 16896
rect 3995 16831 4315 16832
rect 10098 16896 10418 16897
rect 10098 16832 10106 16896
rect 10170 16832 10186 16896
rect 10250 16832 10266 16896
rect 10330 16832 10346 16896
rect 10410 16832 10418 16896
rect 10098 16831 10418 16832
rect 16200 16896 16520 16897
rect 16200 16832 16208 16896
rect 16272 16832 16288 16896
rect 16352 16832 16368 16896
rect 16432 16832 16448 16896
rect 16512 16832 16520 16896
rect 16200 16831 16520 16832
rect 7046 16352 7366 16353
rect 7046 16288 7054 16352
rect 7118 16288 7134 16352
rect 7198 16288 7214 16352
rect 7278 16288 7294 16352
rect 7358 16288 7366 16352
rect 7046 16287 7366 16288
rect 13149 16352 13469 16353
rect 13149 16288 13157 16352
rect 13221 16288 13237 16352
rect 13301 16288 13317 16352
rect 13381 16288 13397 16352
rect 13461 16288 13469 16352
rect 13149 16287 13469 16288
rect 3995 15808 4315 15809
rect 3995 15744 4003 15808
rect 4067 15744 4083 15808
rect 4147 15744 4163 15808
rect 4227 15744 4243 15808
rect 4307 15744 4315 15808
rect 3995 15743 4315 15744
rect 10098 15808 10418 15809
rect 10098 15744 10106 15808
rect 10170 15744 10186 15808
rect 10250 15744 10266 15808
rect 10330 15744 10346 15808
rect 10410 15744 10418 15808
rect 10098 15743 10418 15744
rect 16200 15808 16520 15809
rect 16200 15744 16208 15808
rect 16272 15744 16288 15808
rect 16352 15744 16368 15808
rect 16432 15744 16448 15808
rect 16512 15744 16520 15808
rect 16200 15743 16520 15744
rect 7046 15264 7366 15265
rect 7046 15200 7054 15264
rect 7118 15200 7134 15264
rect 7198 15200 7214 15264
rect 7278 15200 7294 15264
rect 7358 15200 7366 15264
rect 7046 15199 7366 15200
rect 13149 15264 13469 15265
rect 13149 15200 13157 15264
rect 13221 15200 13237 15264
rect 13301 15200 13317 15264
rect 13381 15200 13397 15264
rect 13461 15200 13469 15264
rect 13149 15199 13469 15200
rect 3995 14720 4315 14721
rect 3995 14656 4003 14720
rect 4067 14656 4083 14720
rect 4147 14656 4163 14720
rect 4227 14656 4243 14720
rect 4307 14656 4315 14720
rect 3995 14655 4315 14656
rect 10098 14720 10418 14721
rect 10098 14656 10106 14720
rect 10170 14656 10186 14720
rect 10250 14656 10266 14720
rect 10330 14656 10346 14720
rect 10410 14656 10418 14720
rect 10098 14655 10418 14656
rect 16200 14720 16520 14721
rect 16200 14656 16208 14720
rect 16272 14656 16288 14720
rect 16352 14656 16368 14720
rect 16432 14656 16448 14720
rect 16512 14656 16520 14720
rect 16200 14655 16520 14656
rect 7046 14176 7366 14177
rect 7046 14112 7054 14176
rect 7118 14112 7134 14176
rect 7198 14112 7214 14176
rect 7278 14112 7294 14176
rect 7358 14112 7366 14176
rect 7046 14111 7366 14112
rect 13149 14176 13469 14177
rect 13149 14112 13157 14176
rect 13221 14112 13237 14176
rect 13301 14112 13317 14176
rect 13381 14112 13397 14176
rect 13461 14112 13469 14176
rect 13149 14111 13469 14112
rect 3995 13632 4315 13633
rect 3995 13568 4003 13632
rect 4067 13568 4083 13632
rect 4147 13568 4163 13632
rect 4227 13568 4243 13632
rect 4307 13568 4315 13632
rect 3995 13567 4315 13568
rect 10098 13632 10418 13633
rect 10098 13568 10106 13632
rect 10170 13568 10186 13632
rect 10250 13568 10266 13632
rect 10330 13568 10346 13632
rect 10410 13568 10418 13632
rect 10098 13567 10418 13568
rect 16200 13632 16520 13633
rect 16200 13568 16208 13632
rect 16272 13568 16288 13632
rect 16352 13568 16368 13632
rect 16432 13568 16448 13632
rect 16512 13568 16520 13632
rect 16200 13567 16520 13568
rect 7046 13088 7366 13089
rect 7046 13024 7054 13088
rect 7118 13024 7134 13088
rect 7198 13024 7214 13088
rect 7278 13024 7294 13088
rect 7358 13024 7366 13088
rect 7046 13023 7366 13024
rect 13149 13088 13469 13089
rect 13149 13024 13157 13088
rect 13221 13024 13237 13088
rect 13301 13024 13317 13088
rect 13381 13024 13397 13088
rect 13461 13024 13469 13088
rect 13149 13023 13469 13024
rect 3995 12544 4315 12545
rect 3995 12480 4003 12544
rect 4067 12480 4083 12544
rect 4147 12480 4163 12544
rect 4227 12480 4243 12544
rect 4307 12480 4315 12544
rect 3995 12479 4315 12480
rect 10098 12544 10418 12545
rect 10098 12480 10106 12544
rect 10170 12480 10186 12544
rect 10250 12480 10266 12544
rect 10330 12480 10346 12544
rect 10410 12480 10418 12544
rect 10098 12479 10418 12480
rect 16200 12544 16520 12545
rect 16200 12480 16208 12544
rect 16272 12480 16288 12544
rect 16352 12480 16368 12544
rect 16432 12480 16448 12544
rect 16512 12480 16520 12544
rect 16200 12479 16520 12480
rect 7046 12000 7366 12001
rect 7046 11936 7054 12000
rect 7118 11936 7134 12000
rect 7198 11936 7214 12000
rect 7278 11936 7294 12000
rect 7358 11936 7366 12000
rect 7046 11935 7366 11936
rect 13149 12000 13469 12001
rect 13149 11936 13157 12000
rect 13221 11936 13237 12000
rect 13301 11936 13317 12000
rect 13381 11936 13397 12000
rect 13461 11936 13469 12000
rect 13149 11935 13469 11936
rect 3995 11456 4315 11457
rect 0 11386 800 11416
rect 3995 11392 4003 11456
rect 4067 11392 4083 11456
rect 4147 11392 4163 11456
rect 4227 11392 4243 11456
rect 4307 11392 4315 11456
rect 3995 11391 4315 11392
rect 10098 11456 10418 11457
rect 10098 11392 10106 11456
rect 10170 11392 10186 11456
rect 10250 11392 10266 11456
rect 10330 11392 10346 11456
rect 10410 11392 10418 11456
rect 10098 11391 10418 11392
rect 16200 11456 16520 11457
rect 16200 11392 16208 11456
rect 16272 11392 16288 11456
rect 16352 11392 16368 11456
rect 16432 11392 16448 11456
rect 16512 11392 16520 11456
rect 16200 11391 16520 11392
rect 1577 11386 1643 11389
rect 19717 11386 20517 11416
rect 0 11384 1643 11386
rect 0 11328 1582 11384
rect 1638 11328 1643 11384
rect 0 11326 1643 11328
rect 0 11296 800 11326
rect 1577 11323 1643 11326
rect 16622 11326 20517 11386
rect 15837 11250 15903 11253
rect 16622 11250 16682 11326
rect 19717 11296 20517 11326
rect 15837 11248 16682 11250
rect 15837 11192 15842 11248
rect 15898 11192 16682 11248
rect 15837 11190 16682 11192
rect 15837 11187 15903 11190
rect 7046 10912 7366 10913
rect 7046 10848 7054 10912
rect 7118 10848 7134 10912
rect 7198 10848 7214 10912
rect 7278 10848 7294 10912
rect 7358 10848 7366 10912
rect 7046 10847 7366 10848
rect 13149 10912 13469 10913
rect 13149 10848 13157 10912
rect 13221 10848 13237 10912
rect 13301 10848 13317 10912
rect 13381 10848 13397 10912
rect 13461 10848 13469 10912
rect 13149 10847 13469 10848
rect 3995 10368 4315 10369
rect 3995 10304 4003 10368
rect 4067 10304 4083 10368
rect 4147 10304 4163 10368
rect 4227 10304 4243 10368
rect 4307 10304 4315 10368
rect 3995 10303 4315 10304
rect 10098 10368 10418 10369
rect 10098 10304 10106 10368
rect 10170 10304 10186 10368
rect 10250 10304 10266 10368
rect 10330 10304 10346 10368
rect 10410 10304 10418 10368
rect 10098 10303 10418 10304
rect 16200 10368 16520 10369
rect 16200 10304 16208 10368
rect 16272 10304 16288 10368
rect 16352 10304 16368 10368
rect 16432 10304 16448 10368
rect 16512 10304 16520 10368
rect 16200 10303 16520 10304
rect 7046 9824 7366 9825
rect 7046 9760 7054 9824
rect 7118 9760 7134 9824
rect 7198 9760 7214 9824
rect 7278 9760 7294 9824
rect 7358 9760 7366 9824
rect 7046 9759 7366 9760
rect 13149 9824 13469 9825
rect 13149 9760 13157 9824
rect 13221 9760 13237 9824
rect 13301 9760 13317 9824
rect 13381 9760 13397 9824
rect 13461 9760 13469 9824
rect 13149 9759 13469 9760
rect 3995 9280 4315 9281
rect 3995 9216 4003 9280
rect 4067 9216 4083 9280
rect 4147 9216 4163 9280
rect 4227 9216 4243 9280
rect 4307 9216 4315 9280
rect 3995 9215 4315 9216
rect 10098 9280 10418 9281
rect 10098 9216 10106 9280
rect 10170 9216 10186 9280
rect 10250 9216 10266 9280
rect 10330 9216 10346 9280
rect 10410 9216 10418 9280
rect 10098 9215 10418 9216
rect 16200 9280 16520 9281
rect 16200 9216 16208 9280
rect 16272 9216 16288 9280
rect 16352 9216 16368 9280
rect 16432 9216 16448 9280
rect 16512 9216 16520 9280
rect 16200 9215 16520 9216
rect 7046 8736 7366 8737
rect 7046 8672 7054 8736
rect 7118 8672 7134 8736
rect 7198 8672 7214 8736
rect 7278 8672 7294 8736
rect 7358 8672 7366 8736
rect 7046 8671 7366 8672
rect 13149 8736 13469 8737
rect 13149 8672 13157 8736
rect 13221 8672 13237 8736
rect 13301 8672 13317 8736
rect 13381 8672 13397 8736
rect 13461 8672 13469 8736
rect 13149 8671 13469 8672
rect 3995 8192 4315 8193
rect 3995 8128 4003 8192
rect 4067 8128 4083 8192
rect 4147 8128 4163 8192
rect 4227 8128 4243 8192
rect 4307 8128 4315 8192
rect 3995 8127 4315 8128
rect 10098 8192 10418 8193
rect 10098 8128 10106 8192
rect 10170 8128 10186 8192
rect 10250 8128 10266 8192
rect 10330 8128 10346 8192
rect 10410 8128 10418 8192
rect 10098 8127 10418 8128
rect 16200 8192 16520 8193
rect 16200 8128 16208 8192
rect 16272 8128 16288 8192
rect 16352 8128 16368 8192
rect 16432 8128 16448 8192
rect 16512 8128 16520 8192
rect 16200 8127 16520 8128
rect 7046 7648 7366 7649
rect 7046 7584 7054 7648
rect 7118 7584 7134 7648
rect 7198 7584 7214 7648
rect 7278 7584 7294 7648
rect 7358 7584 7366 7648
rect 7046 7583 7366 7584
rect 13149 7648 13469 7649
rect 13149 7584 13157 7648
rect 13221 7584 13237 7648
rect 13301 7584 13317 7648
rect 13381 7584 13397 7648
rect 13461 7584 13469 7648
rect 13149 7583 13469 7584
rect 3995 7104 4315 7105
rect 3995 7040 4003 7104
rect 4067 7040 4083 7104
rect 4147 7040 4163 7104
rect 4227 7040 4243 7104
rect 4307 7040 4315 7104
rect 3995 7039 4315 7040
rect 10098 7104 10418 7105
rect 10098 7040 10106 7104
rect 10170 7040 10186 7104
rect 10250 7040 10266 7104
rect 10330 7040 10346 7104
rect 10410 7040 10418 7104
rect 10098 7039 10418 7040
rect 16200 7104 16520 7105
rect 16200 7040 16208 7104
rect 16272 7040 16288 7104
rect 16352 7040 16368 7104
rect 16432 7040 16448 7104
rect 16512 7040 16520 7104
rect 16200 7039 16520 7040
rect 7046 6560 7366 6561
rect 7046 6496 7054 6560
rect 7118 6496 7134 6560
rect 7198 6496 7214 6560
rect 7278 6496 7294 6560
rect 7358 6496 7366 6560
rect 7046 6495 7366 6496
rect 13149 6560 13469 6561
rect 13149 6496 13157 6560
rect 13221 6496 13237 6560
rect 13301 6496 13317 6560
rect 13381 6496 13397 6560
rect 13461 6496 13469 6560
rect 13149 6495 13469 6496
rect 3995 6016 4315 6017
rect 3995 5952 4003 6016
rect 4067 5952 4083 6016
rect 4147 5952 4163 6016
rect 4227 5952 4243 6016
rect 4307 5952 4315 6016
rect 3995 5951 4315 5952
rect 10098 6016 10418 6017
rect 10098 5952 10106 6016
rect 10170 5952 10186 6016
rect 10250 5952 10266 6016
rect 10330 5952 10346 6016
rect 10410 5952 10418 6016
rect 10098 5951 10418 5952
rect 16200 6016 16520 6017
rect 16200 5952 16208 6016
rect 16272 5952 16288 6016
rect 16352 5952 16368 6016
rect 16432 5952 16448 6016
rect 16512 5952 16520 6016
rect 16200 5951 16520 5952
rect 7046 5472 7366 5473
rect 7046 5408 7054 5472
rect 7118 5408 7134 5472
rect 7198 5408 7214 5472
rect 7278 5408 7294 5472
rect 7358 5408 7366 5472
rect 7046 5407 7366 5408
rect 13149 5472 13469 5473
rect 13149 5408 13157 5472
rect 13221 5408 13237 5472
rect 13301 5408 13317 5472
rect 13381 5408 13397 5472
rect 13461 5408 13469 5472
rect 13149 5407 13469 5408
rect 3995 4928 4315 4929
rect 3995 4864 4003 4928
rect 4067 4864 4083 4928
rect 4147 4864 4163 4928
rect 4227 4864 4243 4928
rect 4307 4864 4315 4928
rect 3995 4863 4315 4864
rect 10098 4928 10418 4929
rect 10098 4864 10106 4928
rect 10170 4864 10186 4928
rect 10250 4864 10266 4928
rect 10330 4864 10346 4928
rect 10410 4864 10418 4928
rect 10098 4863 10418 4864
rect 16200 4928 16520 4929
rect 16200 4864 16208 4928
rect 16272 4864 16288 4928
rect 16352 4864 16368 4928
rect 16432 4864 16448 4928
rect 16512 4864 16520 4928
rect 16200 4863 16520 4864
rect 7046 4384 7366 4385
rect 7046 4320 7054 4384
rect 7118 4320 7134 4384
rect 7198 4320 7214 4384
rect 7278 4320 7294 4384
rect 7358 4320 7366 4384
rect 7046 4319 7366 4320
rect 13149 4384 13469 4385
rect 13149 4320 13157 4384
rect 13221 4320 13237 4384
rect 13301 4320 13317 4384
rect 13381 4320 13397 4384
rect 13461 4320 13469 4384
rect 13149 4319 13469 4320
rect 3995 3840 4315 3841
rect 3995 3776 4003 3840
rect 4067 3776 4083 3840
rect 4147 3776 4163 3840
rect 4227 3776 4243 3840
rect 4307 3776 4315 3840
rect 3995 3775 4315 3776
rect 10098 3840 10418 3841
rect 10098 3776 10106 3840
rect 10170 3776 10186 3840
rect 10250 3776 10266 3840
rect 10330 3776 10346 3840
rect 10410 3776 10418 3840
rect 10098 3775 10418 3776
rect 16200 3840 16520 3841
rect 16200 3776 16208 3840
rect 16272 3776 16288 3840
rect 16352 3776 16368 3840
rect 16432 3776 16448 3840
rect 16512 3776 16520 3840
rect 16200 3775 16520 3776
rect 7046 3296 7366 3297
rect 7046 3232 7054 3296
rect 7118 3232 7134 3296
rect 7198 3232 7214 3296
rect 7278 3232 7294 3296
rect 7358 3232 7366 3296
rect 7046 3231 7366 3232
rect 13149 3296 13469 3297
rect 13149 3232 13157 3296
rect 13221 3232 13237 3296
rect 13301 3232 13317 3296
rect 13381 3232 13397 3296
rect 13461 3232 13469 3296
rect 13149 3231 13469 3232
rect 3995 2752 4315 2753
rect 3995 2688 4003 2752
rect 4067 2688 4083 2752
rect 4147 2688 4163 2752
rect 4227 2688 4243 2752
rect 4307 2688 4315 2752
rect 3995 2687 4315 2688
rect 10098 2752 10418 2753
rect 10098 2688 10106 2752
rect 10170 2688 10186 2752
rect 10250 2688 10266 2752
rect 10330 2688 10346 2752
rect 10410 2688 10418 2752
rect 10098 2687 10418 2688
rect 16200 2752 16520 2753
rect 16200 2688 16208 2752
rect 16272 2688 16288 2752
rect 16352 2688 16368 2752
rect 16432 2688 16448 2752
rect 16512 2688 16520 2752
rect 16200 2687 16520 2688
rect 7046 2208 7366 2209
rect 7046 2144 7054 2208
rect 7118 2144 7134 2208
rect 7198 2144 7214 2208
rect 7278 2144 7294 2208
rect 7358 2144 7366 2208
rect 7046 2143 7366 2144
rect 13149 2208 13469 2209
rect 13149 2144 13157 2208
rect 13221 2144 13237 2208
rect 13301 2144 13317 2208
rect 13381 2144 13397 2208
rect 13461 2144 13469 2208
rect 13149 2143 13469 2144
<< via3 >>
rect 4003 20156 4067 20160
rect 4003 20100 4007 20156
rect 4007 20100 4063 20156
rect 4063 20100 4067 20156
rect 4003 20096 4067 20100
rect 4083 20156 4147 20160
rect 4083 20100 4087 20156
rect 4087 20100 4143 20156
rect 4143 20100 4147 20156
rect 4083 20096 4147 20100
rect 4163 20156 4227 20160
rect 4163 20100 4167 20156
rect 4167 20100 4223 20156
rect 4223 20100 4227 20156
rect 4163 20096 4227 20100
rect 4243 20156 4307 20160
rect 4243 20100 4247 20156
rect 4247 20100 4303 20156
rect 4303 20100 4307 20156
rect 4243 20096 4307 20100
rect 10106 20156 10170 20160
rect 10106 20100 10110 20156
rect 10110 20100 10166 20156
rect 10166 20100 10170 20156
rect 10106 20096 10170 20100
rect 10186 20156 10250 20160
rect 10186 20100 10190 20156
rect 10190 20100 10246 20156
rect 10246 20100 10250 20156
rect 10186 20096 10250 20100
rect 10266 20156 10330 20160
rect 10266 20100 10270 20156
rect 10270 20100 10326 20156
rect 10326 20100 10330 20156
rect 10266 20096 10330 20100
rect 10346 20156 10410 20160
rect 10346 20100 10350 20156
rect 10350 20100 10406 20156
rect 10406 20100 10410 20156
rect 10346 20096 10410 20100
rect 16208 20156 16272 20160
rect 16208 20100 16212 20156
rect 16212 20100 16268 20156
rect 16268 20100 16272 20156
rect 16208 20096 16272 20100
rect 16288 20156 16352 20160
rect 16288 20100 16292 20156
rect 16292 20100 16348 20156
rect 16348 20100 16352 20156
rect 16288 20096 16352 20100
rect 16368 20156 16432 20160
rect 16368 20100 16372 20156
rect 16372 20100 16428 20156
rect 16428 20100 16432 20156
rect 16368 20096 16432 20100
rect 16448 20156 16512 20160
rect 16448 20100 16452 20156
rect 16452 20100 16508 20156
rect 16508 20100 16512 20156
rect 16448 20096 16512 20100
rect 7054 19612 7118 19616
rect 7054 19556 7058 19612
rect 7058 19556 7114 19612
rect 7114 19556 7118 19612
rect 7054 19552 7118 19556
rect 7134 19612 7198 19616
rect 7134 19556 7138 19612
rect 7138 19556 7194 19612
rect 7194 19556 7198 19612
rect 7134 19552 7198 19556
rect 7214 19612 7278 19616
rect 7214 19556 7218 19612
rect 7218 19556 7274 19612
rect 7274 19556 7278 19612
rect 7214 19552 7278 19556
rect 7294 19612 7358 19616
rect 7294 19556 7298 19612
rect 7298 19556 7354 19612
rect 7354 19556 7358 19612
rect 7294 19552 7358 19556
rect 13157 19612 13221 19616
rect 13157 19556 13161 19612
rect 13161 19556 13217 19612
rect 13217 19556 13221 19612
rect 13157 19552 13221 19556
rect 13237 19612 13301 19616
rect 13237 19556 13241 19612
rect 13241 19556 13297 19612
rect 13297 19556 13301 19612
rect 13237 19552 13301 19556
rect 13317 19612 13381 19616
rect 13317 19556 13321 19612
rect 13321 19556 13377 19612
rect 13377 19556 13381 19612
rect 13317 19552 13381 19556
rect 13397 19612 13461 19616
rect 13397 19556 13401 19612
rect 13401 19556 13457 19612
rect 13457 19556 13461 19612
rect 13397 19552 13461 19556
rect 4003 19068 4067 19072
rect 4003 19012 4007 19068
rect 4007 19012 4063 19068
rect 4063 19012 4067 19068
rect 4003 19008 4067 19012
rect 4083 19068 4147 19072
rect 4083 19012 4087 19068
rect 4087 19012 4143 19068
rect 4143 19012 4147 19068
rect 4083 19008 4147 19012
rect 4163 19068 4227 19072
rect 4163 19012 4167 19068
rect 4167 19012 4223 19068
rect 4223 19012 4227 19068
rect 4163 19008 4227 19012
rect 4243 19068 4307 19072
rect 4243 19012 4247 19068
rect 4247 19012 4303 19068
rect 4303 19012 4307 19068
rect 4243 19008 4307 19012
rect 10106 19068 10170 19072
rect 10106 19012 10110 19068
rect 10110 19012 10166 19068
rect 10166 19012 10170 19068
rect 10106 19008 10170 19012
rect 10186 19068 10250 19072
rect 10186 19012 10190 19068
rect 10190 19012 10246 19068
rect 10246 19012 10250 19068
rect 10186 19008 10250 19012
rect 10266 19068 10330 19072
rect 10266 19012 10270 19068
rect 10270 19012 10326 19068
rect 10326 19012 10330 19068
rect 10266 19008 10330 19012
rect 10346 19068 10410 19072
rect 10346 19012 10350 19068
rect 10350 19012 10406 19068
rect 10406 19012 10410 19068
rect 10346 19008 10410 19012
rect 16208 19068 16272 19072
rect 16208 19012 16212 19068
rect 16212 19012 16268 19068
rect 16268 19012 16272 19068
rect 16208 19008 16272 19012
rect 16288 19068 16352 19072
rect 16288 19012 16292 19068
rect 16292 19012 16348 19068
rect 16348 19012 16352 19068
rect 16288 19008 16352 19012
rect 16368 19068 16432 19072
rect 16368 19012 16372 19068
rect 16372 19012 16428 19068
rect 16428 19012 16432 19068
rect 16368 19008 16432 19012
rect 16448 19068 16512 19072
rect 16448 19012 16452 19068
rect 16452 19012 16508 19068
rect 16508 19012 16512 19068
rect 16448 19008 16512 19012
rect 7054 18524 7118 18528
rect 7054 18468 7058 18524
rect 7058 18468 7114 18524
rect 7114 18468 7118 18524
rect 7054 18464 7118 18468
rect 7134 18524 7198 18528
rect 7134 18468 7138 18524
rect 7138 18468 7194 18524
rect 7194 18468 7198 18524
rect 7134 18464 7198 18468
rect 7214 18524 7278 18528
rect 7214 18468 7218 18524
rect 7218 18468 7274 18524
rect 7274 18468 7278 18524
rect 7214 18464 7278 18468
rect 7294 18524 7358 18528
rect 7294 18468 7298 18524
rect 7298 18468 7354 18524
rect 7354 18468 7358 18524
rect 7294 18464 7358 18468
rect 13157 18524 13221 18528
rect 13157 18468 13161 18524
rect 13161 18468 13217 18524
rect 13217 18468 13221 18524
rect 13157 18464 13221 18468
rect 13237 18524 13301 18528
rect 13237 18468 13241 18524
rect 13241 18468 13297 18524
rect 13297 18468 13301 18524
rect 13237 18464 13301 18468
rect 13317 18524 13381 18528
rect 13317 18468 13321 18524
rect 13321 18468 13377 18524
rect 13377 18468 13381 18524
rect 13317 18464 13381 18468
rect 13397 18524 13461 18528
rect 13397 18468 13401 18524
rect 13401 18468 13457 18524
rect 13457 18468 13461 18524
rect 13397 18464 13461 18468
rect 4003 17980 4067 17984
rect 4003 17924 4007 17980
rect 4007 17924 4063 17980
rect 4063 17924 4067 17980
rect 4003 17920 4067 17924
rect 4083 17980 4147 17984
rect 4083 17924 4087 17980
rect 4087 17924 4143 17980
rect 4143 17924 4147 17980
rect 4083 17920 4147 17924
rect 4163 17980 4227 17984
rect 4163 17924 4167 17980
rect 4167 17924 4223 17980
rect 4223 17924 4227 17980
rect 4163 17920 4227 17924
rect 4243 17980 4307 17984
rect 4243 17924 4247 17980
rect 4247 17924 4303 17980
rect 4303 17924 4307 17980
rect 4243 17920 4307 17924
rect 10106 17980 10170 17984
rect 10106 17924 10110 17980
rect 10110 17924 10166 17980
rect 10166 17924 10170 17980
rect 10106 17920 10170 17924
rect 10186 17980 10250 17984
rect 10186 17924 10190 17980
rect 10190 17924 10246 17980
rect 10246 17924 10250 17980
rect 10186 17920 10250 17924
rect 10266 17980 10330 17984
rect 10266 17924 10270 17980
rect 10270 17924 10326 17980
rect 10326 17924 10330 17980
rect 10266 17920 10330 17924
rect 10346 17980 10410 17984
rect 10346 17924 10350 17980
rect 10350 17924 10406 17980
rect 10406 17924 10410 17980
rect 10346 17920 10410 17924
rect 16208 17980 16272 17984
rect 16208 17924 16212 17980
rect 16212 17924 16268 17980
rect 16268 17924 16272 17980
rect 16208 17920 16272 17924
rect 16288 17980 16352 17984
rect 16288 17924 16292 17980
rect 16292 17924 16348 17980
rect 16348 17924 16352 17980
rect 16288 17920 16352 17924
rect 16368 17980 16432 17984
rect 16368 17924 16372 17980
rect 16372 17924 16428 17980
rect 16428 17924 16432 17980
rect 16368 17920 16432 17924
rect 16448 17980 16512 17984
rect 16448 17924 16452 17980
rect 16452 17924 16508 17980
rect 16508 17924 16512 17980
rect 16448 17920 16512 17924
rect 7054 17436 7118 17440
rect 7054 17380 7058 17436
rect 7058 17380 7114 17436
rect 7114 17380 7118 17436
rect 7054 17376 7118 17380
rect 7134 17436 7198 17440
rect 7134 17380 7138 17436
rect 7138 17380 7194 17436
rect 7194 17380 7198 17436
rect 7134 17376 7198 17380
rect 7214 17436 7278 17440
rect 7214 17380 7218 17436
rect 7218 17380 7274 17436
rect 7274 17380 7278 17436
rect 7214 17376 7278 17380
rect 7294 17436 7358 17440
rect 7294 17380 7298 17436
rect 7298 17380 7354 17436
rect 7354 17380 7358 17436
rect 7294 17376 7358 17380
rect 13157 17436 13221 17440
rect 13157 17380 13161 17436
rect 13161 17380 13217 17436
rect 13217 17380 13221 17436
rect 13157 17376 13221 17380
rect 13237 17436 13301 17440
rect 13237 17380 13241 17436
rect 13241 17380 13297 17436
rect 13297 17380 13301 17436
rect 13237 17376 13301 17380
rect 13317 17436 13381 17440
rect 13317 17380 13321 17436
rect 13321 17380 13377 17436
rect 13377 17380 13381 17436
rect 13317 17376 13381 17380
rect 13397 17436 13461 17440
rect 13397 17380 13401 17436
rect 13401 17380 13457 17436
rect 13457 17380 13461 17436
rect 13397 17376 13461 17380
rect 4003 16892 4067 16896
rect 4003 16836 4007 16892
rect 4007 16836 4063 16892
rect 4063 16836 4067 16892
rect 4003 16832 4067 16836
rect 4083 16892 4147 16896
rect 4083 16836 4087 16892
rect 4087 16836 4143 16892
rect 4143 16836 4147 16892
rect 4083 16832 4147 16836
rect 4163 16892 4227 16896
rect 4163 16836 4167 16892
rect 4167 16836 4223 16892
rect 4223 16836 4227 16892
rect 4163 16832 4227 16836
rect 4243 16892 4307 16896
rect 4243 16836 4247 16892
rect 4247 16836 4303 16892
rect 4303 16836 4307 16892
rect 4243 16832 4307 16836
rect 10106 16892 10170 16896
rect 10106 16836 10110 16892
rect 10110 16836 10166 16892
rect 10166 16836 10170 16892
rect 10106 16832 10170 16836
rect 10186 16892 10250 16896
rect 10186 16836 10190 16892
rect 10190 16836 10246 16892
rect 10246 16836 10250 16892
rect 10186 16832 10250 16836
rect 10266 16892 10330 16896
rect 10266 16836 10270 16892
rect 10270 16836 10326 16892
rect 10326 16836 10330 16892
rect 10266 16832 10330 16836
rect 10346 16892 10410 16896
rect 10346 16836 10350 16892
rect 10350 16836 10406 16892
rect 10406 16836 10410 16892
rect 10346 16832 10410 16836
rect 16208 16892 16272 16896
rect 16208 16836 16212 16892
rect 16212 16836 16268 16892
rect 16268 16836 16272 16892
rect 16208 16832 16272 16836
rect 16288 16892 16352 16896
rect 16288 16836 16292 16892
rect 16292 16836 16348 16892
rect 16348 16836 16352 16892
rect 16288 16832 16352 16836
rect 16368 16892 16432 16896
rect 16368 16836 16372 16892
rect 16372 16836 16428 16892
rect 16428 16836 16432 16892
rect 16368 16832 16432 16836
rect 16448 16892 16512 16896
rect 16448 16836 16452 16892
rect 16452 16836 16508 16892
rect 16508 16836 16512 16892
rect 16448 16832 16512 16836
rect 7054 16348 7118 16352
rect 7054 16292 7058 16348
rect 7058 16292 7114 16348
rect 7114 16292 7118 16348
rect 7054 16288 7118 16292
rect 7134 16348 7198 16352
rect 7134 16292 7138 16348
rect 7138 16292 7194 16348
rect 7194 16292 7198 16348
rect 7134 16288 7198 16292
rect 7214 16348 7278 16352
rect 7214 16292 7218 16348
rect 7218 16292 7274 16348
rect 7274 16292 7278 16348
rect 7214 16288 7278 16292
rect 7294 16348 7358 16352
rect 7294 16292 7298 16348
rect 7298 16292 7354 16348
rect 7354 16292 7358 16348
rect 7294 16288 7358 16292
rect 13157 16348 13221 16352
rect 13157 16292 13161 16348
rect 13161 16292 13217 16348
rect 13217 16292 13221 16348
rect 13157 16288 13221 16292
rect 13237 16348 13301 16352
rect 13237 16292 13241 16348
rect 13241 16292 13297 16348
rect 13297 16292 13301 16348
rect 13237 16288 13301 16292
rect 13317 16348 13381 16352
rect 13317 16292 13321 16348
rect 13321 16292 13377 16348
rect 13377 16292 13381 16348
rect 13317 16288 13381 16292
rect 13397 16348 13461 16352
rect 13397 16292 13401 16348
rect 13401 16292 13457 16348
rect 13457 16292 13461 16348
rect 13397 16288 13461 16292
rect 4003 15804 4067 15808
rect 4003 15748 4007 15804
rect 4007 15748 4063 15804
rect 4063 15748 4067 15804
rect 4003 15744 4067 15748
rect 4083 15804 4147 15808
rect 4083 15748 4087 15804
rect 4087 15748 4143 15804
rect 4143 15748 4147 15804
rect 4083 15744 4147 15748
rect 4163 15804 4227 15808
rect 4163 15748 4167 15804
rect 4167 15748 4223 15804
rect 4223 15748 4227 15804
rect 4163 15744 4227 15748
rect 4243 15804 4307 15808
rect 4243 15748 4247 15804
rect 4247 15748 4303 15804
rect 4303 15748 4307 15804
rect 4243 15744 4307 15748
rect 10106 15804 10170 15808
rect 10106 15748 10110 15804
rect 10110 15748 10166 15804
rect 10166 15748 10170 15804
rect 10106 15744 10170 15748
rect 10186 15804 10250 15808
rect 10186 15748 10190 15804
rect 10190 15748 10246 15804
rect 10246 15748 10250 15804
rect 10186 15744 10250 15748
rect 10266 15804 10330 15808
rect 10266 15748 10270 15804
rect 10270 15748 10326 15804
rect 10326 15748 10330 15804
rect 10266 15744 10330 15748
rect 10346 15804 10410 15808
rect 10346 15748 10350 15804
rect 10350 15748 10406 15804
rect 10406 15748 10410 15804
rect 10346 15744 10410 15748
rect 16208 15804 16272 15808
rect 16208 15748 16212 15804
rect 16212 15748 16268 15804
rect 16268 15748 16272 15804
rect 16208 15744 16272 15748
rect 16288 15804 16352 15808
rect 16288 15748 16292 15804
rect 16292 15748 16348 15804
rect 16348 15748 16352 15804
rect 16288 15744 16352 15748
rect 16368 15804 16432 15808
rect 16368 15748 16372 15804
rect 16372 15748 16428 15804
rect 16428 15748 16432 15804
rect 16368 15744 16432 15748
rect 16448 15804 16512 15808
rect 16448 15748 16452 15804
rect 16452 15748 16508 15804
rect 16508 15748 16512 15804
rect 16448 15744 16512 15748
rect 7054 15260 7118 15264
rect 7054 15204 7058 15260
rect 7058 15204 7114 15260
rect 7114 15204 7118 15260
rect 7054 15200 7118 15204
rect 7134 15260 7198 15264
rect 7134 15204 7138 15260
rect 7138 15204 7194 15260
rect 7194 15204 7198 15260
rect 7134 15200 7198 15204
rect 7214 15260 7278 15264
rect 7214 15204 7218 15260
rect 7218 15204 7274 15260
rect 7274 15204 7278 15260
rect 7214 15200 7278 15204
rect 7294 15260 7358 15264
rect 7294 15204 7298 15260
rect 7298 15204 7354 15260
rect 7354 15204 7358 15260
rect 7294 15200 7358 15204
rect 13157 15260 13221 15264
rect 13157 15204 13161 15260
rect 13161 15204 13217 15260
rect 13217 15204 13221 15260
rect 13157 15200 13221 15204
rect 13237 15260 13301 15264
rect 13237 15204 13241 15260
rect 13241 15204 13297 15260
rect 13297 15204 13301 15260
rect 13237 15200 13301 15204
rect 13317 15260 13381 15264
rect 13317 15204 13321 15260
rect 13321 15204 13377 15260
rect 13377 15204 13381 15260
rect 13317 15200 13381 15204
rect 13397 15260 13461 15264
rect 13397 15204 13401 15260
rect 13401 15204 13457 15260
rect 13457 15204 13461 15260
rect 13397 15200 13461 15204
rect 4003 14716 4067 14720
rect 4003 14660 4007 14716
rect 4007 14660 4063 14716
rect 4063 14660 4067 14716
rect 4003 14656 4067 14660
rect 4083 14716 4147 14720
rect 4083 14660 4087 14716
rect 4087 14660 4143 14716
rect 4143 14660 4147 14716
rect 4083 14656 4147 14660
rect 4163 14716 4227 14720
rect 4163 14660 4167 14716
rect 4167 14660 4223 14716
rect 4223 14660 4227 14716
rect 4163 14656 4227 14660
rect 4243 14716 4307 14720
rect 4243 14660 4247 14716
rect 4247 14660 4303 14716
rect 4303 14660 4307 14716
rect 4243 14656 4307 14660
rect 10106 14716 10170 14720
rect 10106 14660 10110 14716
rect 10110 14660 10166 14716
rect 10166 14660 10170 14716
rect 10106 14656 10170 14660
rect 10186 14716 10250 14720
rect 10186 14660 10190 14716
rect 10190 14660 10246 14716
rect 10246 14660 10250 14716
rect 10186 14656 10250 14660
rect 10266 14716 10330 14720
rect 10266 14660 10270 14716
rect 10270 14660 10326 14716
rect 10326 14660 10330 14716
rect 10266 14656 10330 14660
rect 10346 14716 10410 14720
rect 10346 14660 10350 14716
rect 10350 14660 10406 14716
rect 10406 14660 10410 14716
rect 10346 14656 10410 14660
rect 16208 14716 16272 14720
rect 16208 14660 16212 14716
rect 16212 14660 16268 14716
rect 16268 14660 16272 14716
rect 16208 14656 16272 14660
rect 16288 14716 16352 14720
rect 16288 14660 16292 14716
rect 16292 14660 16348 14716
rect 16348 14660 16352 14716
rect 16288 14656 16352 14660
rect 16368 14716 16432 14720
rect 16368 14660 16372 14716
rect 16372 14660 16428 14716
rect 16428 14660 16432 14716
rect 16368 14656 16432 14660
rect 16448 14716 16512 14720
rect 16448 14660 16452 14716
rect 16452 14660 16508 14716
rect 16508 14660 16512 14716
rect 16448 14656 16512 14660
rect 7054 14172 7118 14176
rect 7054 14116 7058 14172
rect 7058 14116 7114 14172
rect 7114 14116 7118 14172
rect 7054 14112 7118 14116
rect 7134 14172 7198 14176
rect 7134 14116 7138 14172
rect 7138 14116 7194 14172
rect 7194 14116 7198 14172
rect 7134 14112 7198 14116
rect 7214 14172 7278 14176
rect 7214 14116 7218 14172
rect 7218 14116 7274 14172
rect 7274 14116 7278 14172
rect 7214 14112 7278 14116
rect 7294 14172 7358 14176
rect 7294 14116 7298 14172
rect 7298 14116 7354 14172
rect 7354 14116 7358 14172
rect 7294 14112 7358 14116
rect 13157 14172 13221 14176
rect 13157 14116 13161 14172
rect 13161 14116 13217 14172
rect 13217 14116 13221 14172
rect 13157 14112 13221 14116
rect 13237 14172 13301 14176
rect 13237 14116 13241 14172
rect 13241 14116 13297 14172
rect 13297 14116 13301 14172
rect 13237 14112 13301 14116
rect 13317 14172 13381 14176
rect 13317 14116 13321 14172
rect 13321 14116 13377 14172
rect 13377 14116 13381 14172
rect 13317 14112 13381 14116
rect 13397 14172 13461 14176
rect 13397 14116 13401 14172
rect 13401 14116 13457 14172
rect 13457 14116 13461 14172
rect 13397 14112 13461 14116
rect 4003 13628 4067 13632
rect 4003 13572 4007 13628
rect 4007 13572 4063 13628
rect 4063 13572 4067 13628
rect 4003 13568 4067 13572
rect 4083 13628 4147 13632
rect 4083 13572 4087 13628
rect 4087 13572 4143 13628
rect 4143 13572 4147 13628
rect 4083 13568 4147 13572
rect 4163 13628 4227 13632
rect 4163 13572 4167 13628
rect 4167 13572 4223 13628
rect 4223 13572 4227 13628
rect 4163 13568 4227 13572
rect 4243 13628 4307 13632
rect 4243 13572 4247 13628
rect 4247 13572 4303 13628
rect 4303 13572 4307 13628
rect 4243 13568 4307 13572
rect 10106 13628 10170 13632
rect 10106 13572 10110 13628
rect 10110 13572 10166 13628
rect 10166 13572 10170 13628
rect 10106 13568 10170 13572
rect 10186 13628 10250 13632
rect 10186 13572 10190 13628
rect 10190 13572 10246 13628
rect 10246 13572 10250 13628
rect 10186 13568 10250 13572
rect 10266 13628 10330 13632
rect 10266 13572 10270 13628
rect 10270 13572 10326 13628
rect 10326 13572 10330 13628
rect 10266 13568 10330 13572
rect 10346 13628 10410 13632
rect 10346 13572 10350 13628
rect 10350 13572 10406 13628
rect 10406 13572 10410 13628
rect 10346 13568 10410 13572
rect 16208 13628 16272 13632
rect 16208 13572 16212 13628
rect 16212 13572 16268 13628
rect 16268 13572 16272 13628
rect 16208 13568 16272 13572
rect 16288 13628 16352 13632
rect 16288 13572 16292 13628
rect 16292 13572 16348 13628
rect 16348 13572 16352 13628
rect 16288 13568 16352 13572
rect 16368 13628 16432 13632
rect 16368 13572 16372 13628
rect 16372 13572 16428 13628
rect 16428 13572 16432 13628
rect 16368 13568 16432 13572
rect 16448 13628 16512 13632
rect 16448 13572 16452 13628
rect 16452 13572 16508 13628
rect 16508 13572 16512 13628
rect 16448 13568 16512 13572
rect 7054 13084 7118 13088
rect 7054 13028 7058 13084
rect 7058 13028 7114 13084
rect 7114 13028 7118 13084
rect 7054 13024 7118 13028
rect 7134 13084 7198 13088
rect 7134 13028 7138 13084
rect 7138 13028 7194 13084
rect 7194 13028 7198 13084
rect 7134 13024 7198 13028
rect 7214 13084 7278 13088
rect 7214 13028 7218 13084
rect 7218 13028 7274 13084
rect 7274 13028 7278 13084
rect 7214 13024 7278 13028
rect 7294 13084 7358 13088
rect 7294 13028 7298 13084
rect 7298 13028 7354 13084
rect 7354 13028 7358 13084
rect 7294 13024 7358 13028
rect 13157 13084 13221 13088
rect 13157 13028 13161 13084
rect 13161 13028 13217 13084
rect 13217 13028 13221 13084
rect 13157 13024 13221 13028
rect 13237 13084 13301 13088
rect 13237 13028 13241 13084
rect 13241 13028 13297 13084
rect 13297 13028 13301 13084
rect 13237 13024 13301 13028
rect 13317 13084 13381 13088
rect 13317 13028 13321 13084
rect 13321 13028 13377 13084
rect 13377 13028 13381 13084
rect 13317 13024 13381 13028
rect 13397 13084 13461 13088
rect 13397 13028 13401 13084
rect 13401 13028 13457 13084
rect 13457 13028 13461 13084
rect 13397 13024 13461 13028
rect 4003 12540 4067 12544
rect 4003 12484 4007 12540
rect 4007 12484 4063 12540
rect 4063 12484 4067 12540
rect 4003 12480 4067 12484
rect 4083 12540 4147 12544
rect 4083 12484 4087 12540
rect 4087 12484 4143 12540
rect 4143 12484 4147 12540
rect 4083 12480 4147 12484
rect 4163 12540 4227 12544
rect 4163 12484 4167 12540
rect 4167 12484 4223 12540
rect 4223 12484 4227 12540
rect 4163 12480 4227 12484
rect 4243 12540 4307 12544
rect 4243 12484 4247 12540
rect 4247 12484 4303 12540
rect 4303 12484 4307 12540
rect 4243 12480 4307 12484
rect 10106 12540 10170 12544
rect 10106 12484 10110 12540
rect 10110 12484 10166 12540
rect 10166 12484 10170 12540
rect 10106 12480 10170 12484
rect 10186 12540 10250 12544
rect 10186 12484 10190 12540
rect 10190 12484 10246 12540
rect 10246 12484 10250 12540
rect 10186 12480 10250 12484
rect 10266 12540 10330 12544
rect 10266 12484 10270 12540
rect 10270 12484 10326 12540
rect 10326 12484 10330 12540
rect 10266 12480 10330 12484
rect 10346 12540 10410 12544
rect 10346 12484 10350 12540
rect 10350 12484 10406 12540
rect 10406 12484 10410 12540
rect 10346 12480 10410 12484
rect 16208 12540 16272 12544
rect 16208 12484 16212 12540
rect 16212 12484 16268 12540
rect 16268 12484 16272 12540
rect 16208 12480 16272 12484
rect 16288 12540 16352 12544
rect 16288 12484 16292 12540
rect 16292 12484 16348 12540
rect 16348 12484 16352 12540
rect 16288 12480 16352 12484
rect 16368 12540 16432 12544
rect 16368 12484 16372 12540
rect 16372 12484 16428 12540
rect 16428 12484 16432 12540
rect 16368 12480 16432 12484
rect 16448 12540 16512 12544
rect 16448 12484 16452 12540
rect 16452 12484 16508 12540
rect 16508 12484 16512 12540
rect 16448 12480 16512 12484
rect 7054 11996 7118 12000
rect 7054 11940 7058 11996
rect 7058 11940 7114 11996
rect 7114 11940 7118 11996
rect 7054 11936 7118 11940
rect 7134 11996 7198 12000
rect 7134 11940 7138 11996
rect 7138 11940 7194 11996
rect 7194 11940 7198 11996
rect 7134 11936 7198 11940
rect 7214 11996 7278 12000
rect 7214 11940 7218 11996
rect 7218 11940 7274 11996
rect 7274 11940 7278 11996
rect 7214 11936 7278 11940
rect 7294 11996 7358 12000
rect 7294 11940 7298 11996
rect 7298 11940 7354 11996
rect 7354 11940 7358 11996
rect 7294 11936 7358 11940
rect 13157 11996 13221 12000
rect 13157 11940 13161 11996
rect 13161 11940 13217 11996
rect 13217 11940 13221 11996
rect 13157 11936 13221 11940
rect 13237 11996 13301 12000
rect 13237 11940 13241 11996
rect 13241 11940 13297 11996
rect 13297 11940 13301 11996
rect 13237 11936 13301 11940
rect 13317 11996 13381 12000
rect 13317 11940 13321 11996
rect 13321 11940 13377 11996
rect 13377 11940 13381 11996
rect 13317 11936 13381 11940
rect 13397 11996 13461 12000
rect 13397 11940 13401 11996
rect 13401 11940 13457 11996
rect 13457 11940 13461 11996
rect 13397 11936 13461 11940
rect 4003 11452 4067 11456
rect 4003 11396 4007 11452
rect 4007 11396 4063 11452
rect 4063 11396 4067 11452
rect 4003 11392 4067 11396
rect 4083 11452 4147 11456
rect 4083 11396 4087 11452
rect 4087 11396 4143 11452
rect 4143 11396 4147 11452
rect 4083 11392 4147 11396
rect 4163 11452 4227 11456
rect 4163 11396 4167 11452
rect 4167 11396 4223 11452
rect 4223 11396 4227 11452
rect 4163 11392 4227 11396
rect 4243 11452 4307 11456
rect 4243 11396 4247 11452
rect 4247 11396 4303 11452
rect 4303 11396 4307 11452
rect 4243 11392 4307 11396
rect 10106 11452 10170 11456
rect 10106 11396 10110 11452
rect 10110 11396 10166 11452
rect 10166 11396 10170 11452
rect 10106 11392 10170 11396
rect 10186 11452 10250 11456
rect 10186 11396 10190 11452
rect 10190 11396 10246 11452
rect 10246 11396 10250 11452
rect 10186 11392 10250 11396
rect 10266 11452 10330 11456
rect 10266 11396 10270 11452
rect 10270 11396 10326 11452
rect 10326 11396 10330 11452
rect 10266 11392 10330 11396
rect 10346 11452 10410 11456
rect 10346 11396 10350 11452
rect 10350 11396 10406 11452
rect 10406 11396 10410 11452
rect 10346 11392 10410 11396
rect 16208 11452 16272 11456
rect 16208 11396 16212 11452
rect 16212 11396 16268 11452
rect 16268 11396 16272 11452
rect 16208 11392 16272 11396
rect 16288 11452 16352 11456
rect 16288 11396 16292 11452
rect 16292 11396 16348 11452
rect 16348 11396 16352 11452
rect 16288 11392 16352 11396
rect 16368 11452 16432 11456
rect 16368 11396 16372 11452
rect 16372 11396 16428 11452
rect 16428 11396 16432 11452
rect 16368 11392 16432 11396
rect 16448 11452 16512 11456
rect 16448 11396 16452 11452
rect 16452 11396 16508 11452
rect 16508 11396 16512 11452
rect 16448 11392 16512 11396
rect 7054 10908 7118 10912
rect 7054 10852 7058 10908
rect 7058 10852 7114 10908
rect 7114 10852 7118 10908
rect 7054 10848 7118 10852
rect 7134 10908 7198 10912
rect 7134 10852 7138 10908
rect 7138 10852 7194 10908
rect 7194 10852 7198 10908
rect 7134 10848 7198 10852
rect 7214 10908 7278 10912
rect 7214 10852 7218 10908
rect 7218 10852 7274 10908
rect 7274 10852 7278 10908
rect 7214 10848 7278 10852
rect 7294 10908 7358 10912
rect 7294 10852 7298 10908
rect 7298 10852 7354 10908
rect 7354 10852 7358 10908
rect 7294 10848 7358 10852
rect 13157 10908 13221 10912
rect 13157 10852 13161 10908
rect 13161 10852 13217 10908
rect 13217 10852 13221 10908
rect 13157 10848 13221 10852
rect 13237 10908 13301 10912
rect 13237 10852 13241 10908
rect 13241 10852 13297 10908
rect 13297 10852 13301 10908
rect 13237 10848 13301 10852
rect 13317 10908 13381 10912
rect 13317 10852 13321 10908
rect 13321 10852 13377 10908
rect 13377 10852 13381 10908
rect 13317 10848 13381 10852
rect 13397 10908 13461 10912
rect 13397 10852 13401 10908
rect 13401 10852 13457 10908
rect 13457 10852 13461 10908
rect 13397 10848 13461 10852
rect 4003 10364 4067 10368
rect 4003 10308 4007 10364
rect 4007 10308 4063 10364
rect 4063 10308 4067 10364
rect 4003 10304 4067 10308
rect 4083 10364 4147 10368
rect 4083 10308 4087 10364
rect 4087 10308 4143 10364
rect 4143 10308 4147 10364
rect 4083 10304 4147 10308
rect 4163 10364 4227 10368
rect 4163 10308 4167 10364
rect 4167 10308 4223 10364
rect 4223 10308 4227 10364
rect 4163 10304 4227 10308
rect 4243 10364 4307 10368
rect 4243 10308 4247 10364
rect 4247 10308 4303 10364
rect 4303 10308 4307 10364
rect 4243 10304 4307 10308
rect 10106 10364 10170 10368
rect 10106 10308 10110 10364
rect 10110 10308 10166 10364
rect 10166 10308 10170 10364
rect 10106 10304 10170 10308
rect 10186 10364 10250 10368
rect 10186 10308 10190 10364
rect 10190 10308 10246 10364
rect 10246 10308 10250 10364
rect 10186 10304 10250 10308
rect 10266 10364 10330 10368
rect 10266 10308 10270 10364
rect 10270 10308 10326 10364
rect 10326 10308 10330 10364
rect 10266 10304 10330 10308
rect 10346 10364 10410 10368
rect 10346 10308 10350 10364
rect 10350 10308 10406 10364
rect 10406 10308 10410 10364
rect 10346 10304 10410 10308
rect 16208 10364 16272 10368
rect 16208 10308 16212 10364
rect 16212 10308 16268 10364
rect 16268 10308 16272 10364
rect 16208 10304 16272 10308
rect 16288 10364 16352 10368
rect 16288 10308 16292 10364
rect 16292 10308 16348 10364
rect 16348 10308 16352 10364
rect 16288 10304 16352 10308
rect 16368 10364 16432 10368
rect 16368 10308 16372 10364
rect 16372 10308 16428 10364
rect 16428 10308 16432 10364
rect 16368 10304 16432 10308
rect 16448 10364 16512 10368
rect 16448 10308 16452 10364
rect 16452 10308 16508 10364
rect 16508 10308 16512 10364
rect 16448 10304 16512 10308
rect 7054 9820 7118 9824
rect 7054 9764 7058 9820
rect 7058 9764 7114 9820
rect 7114 9764 7118 9820
rect 7054 9760 7118 9764
rect 7134 9820 7198 9824
rect 7134 9764 7138 9820
rect 7138 9764 7194 9820
rect 7194 9764 7198 9820
rect 7134 9760 7198 9764
rect 7214 9820 7278 9824
rect 7214 9764 7218 9820
rect 7218 9764 7274 9820
rect 7274 9764 7278 9820
rect 7214 9760 7278 9764
rect 7294 9820 7358 9824
rect 7294 9764 7298 9820
rect 7298 9764 7354 9820
rect 7354 9764 7358 9820
rect 7294 9760 7358 9764
rect 13157 9820 13221 9824
rect 13157 9764 13161 9820
rect 13161 9764 13217 9820
rect 13217 9764 13221 9820
rect 13157 9760 13221 9764
rect 13237 9820 13301 9824
rect 13237 9764 13241 9820
rect 13241 9764 13297 9820
rect 13297 9764 13301 9820
rect 13237 9760 13301 9764
rect 13317 9820 13381 9824
rect 13317 9764 13321 9820
rect 13321 9764 13377 9820
rect 13377 9764 13381 9820
rect 13317 9760 13381 9764
rect 13397 9820 13461 9824
rect 13397 9764 13401 9820
rect 13401 9764 13457 9820
rect 13457 9764 13461 9820
rect 13397 9760 13461 9764
rect 4003 9276 4067 9280
rect 4003 9220 4007 9276
rect 4007 9220 4063 9276
rect 4063 9220 4067 9276
rect 4003 9216 4067 9220
rect 4083 9276 4147 9280
rect 4083 9220 4087 9276
rect 4087 9220 4143 9276
rect 4143 9220 4147 9276
rect 4083 9216 4147 9220
rect 4163 9276 4227 9280
rect 4163 9220 4167 9276
rect 4167 9220 4223 9276
rect 4223 9220 4227 9276
rect 4163 9216 4227 9220
rect 4243 9276 4307 9280
rect 4243 9220 4247 9276
rect 4247 9220 4303 9276
rect 4303 9220 4307 9276
rect 4243 9216 4307 9220
rect 10106 9276 10170 9280
rect 10106 9220 10110 9276
rect 10110 9220 10166 9276
rect 10166 9220 10170 9276
rect 10106 9216 10170 9220
rect 10186 9276 10250 9280
rect 10186 9220 10190 9276
rect 10190 9220 10246 9276
rect 10246 9220 10250 9276
rect 10186 9216 10250 9220
rect 10266 9276 10330 9280
rect 10266 9220 10270 9276
rect 10270 9220 10326 9276
rect 10326 9220 10330 9276
rect 10266 9216 10330 9220
rect 10346 9276 10410 9280
rect 10346 9220 10350 9276
rect 10350 9220 10406 9276
rect 10406 9220 10410 9276
rect 10346 9216 10410 9220
rect 16208 9276 16272 9280
rect 16208 9220 16212 9276
rect 16212 9220 16268 9276
rect 16268 9220 16272 9276
rect 16208 9216 16272 9220
rect 16288 9276 16352 9280
rect 16288 9220 16292 9276
rect 16292 9220 16348 9276
rect 16348 9220 16352 9276
rect 16288 9216 16352 9220
rect 16368 9276 16432 9280
rect 16368 9220 16372 9276
rect 16372 9220 16428 9276
rect 16428 9220 16432 9276
rect 16368 9216 16432 9220
rect 16448 9276 16512 9280
rect 16448 9220 16452 9276
rect 16452 9220 16508 9276
rect 16508 9220 16512 9276
rect 16448 9216 16512 9220
rect 7054 8732 7118 8736
rect 7054 8676 7058 8732
rect 7058 8676 7114 8732
rect 7114 8676 7118 8732
rect 7054 8672 7118 8676
rect 7134 8732 7198 8736
rect 7134 8676 7138 8732
rect 7138 8676 7194 8732
rect 7194 8676 7198 8732
rect 7134 8672 7198 8676
rect 7214 8732 7278 8736
rect 7214 8676 7218 8732
rect 7218 8676 7274 8732
rect 7274 8676 7278 8732
rect 7214 8672 7278 8676
rect 7294 8732 7358 8736
rect 7294 8676 7298 8732
rect 7298 8676 7354 8732
rect 7354 8676 7358 8732
rect 7294 8672 7358 8676
rect 13157 8732 13221 8736
rect 13157 8676 13161 8732
rect 13161 8676 13217 8732
rect 13217 8676 13221 8732
rect 13157 8672 13221 8676
rect 13237 8732 13301 8736
rect 13237 8676 13241 8732
rect 13241 8676 13297 8732
rect 13297 8676 13301 8732
rect 13237 8672 13301 8676
rect 13317 8732 13381 8736
rect 13317 8676 13321 8732
rect 13321 8676 13377 8732
rect 13377 8676 13381 8732
rect 13317 8672 13381 8676
rect 13397 8732 13461 8736
rect 13397 8676 13401 8732
rect 13401 8676 13457 8732
rect 13457 8676 13461 8732
rect 13397 8672 13461 8676
rect 4003 8188 4067 8192
rect 4003 8132 4007 8188
rect 4007 8132 4063 8188
rect 4063 8132 4067 8188
rect 4003 8128 4067 8132
rect 4083 8188 4147 8192
rect 4083 8132 4087 8188
rect 4087 8132 4143 8188
rect 4143 8132 4147 8188
rect 4083 8128 4147 8132
rect 4163 8188 4227 8192
rect 4163 8132 4167 8188
rect 4167 8132 4223 8188
rect 4223 8132 4227 8188
rect 4163 8128 4227 8132
rect 4243 8188 4307 8192
rect 4243 8132 4247 8188
rect 4247 8132 4303 8188
rect 4303 8132 4307 8188
rect 4243 8128 4307 8132
rect 10106 8188 10170 8192
rect 10106 8132 10110 8188
rect 10110 8132 10166 8188
rect 10166 8132 10170 8188
rect 10106 8128 10170 8132
rect 10186 8188 10250 8192
rect 10186 8132 10190 8188
rect 10190 8132 10246 8188
rect 10246 8132 10250 8188
rect 10186 8128 10250 8132
rect 10266 8188 10330 8192
rect 10266 8132 10270 8188
rect 10270 8132 10326 8188
rect 10326 8132 10330 8188
rect 10266 8128 10330 8132
rect 10346 8188 10410 8192
rect 10346 8132 10350 8188
rect 10350 8132 10406 8188
rect 10406 8132 10410 8188
rect 10346 8128 10410 8132
rect 16208 8188 16272 8192
rect 16208 8132 16212 8188
rect 16212 8132 16268 8188
rect 16268 8132 16272 8188
rect 16208 8128 16272 8132
rect 16288 8188 16352 8192
rect 16288 8132 16292 8188
rect 16292 8132 16348 8188
rect 16348 8132 16352 8188
rect 16288 8128 16352 8132
rect 16368 8188 16432 8192
rect 16368 8132 16372 8188
rect 16372 8132 16428 8188
rect 16428 8132 16432 8188
rect 16368 8128 16432 8132
rect 16448 8188 16512 8192
rect 16448 8132 16452 8188
rect 16452 8132 16508 8188
rect 16508 8132 16512 8188
rect 16448 8128 16512 8132
rect 7054 7644 7118 7648
rect 7054 7588 7058 7644
rect 7058 7588 7114 7644
rect 7114 7588 7118 7644
rect 7054 7584 7118 7588
rect 7134 7644 7198 7648
rect 7134 7588 7138 7644
rect 7138 7588 7194 7644
rect 7194 7588 7198 7644
rect 7134 7584 7198 7588
rect 7214 7644 7278 7648
rect 7214 7588 7218 7644
rect 7218 7588 7274 7644
rect 7274 7588 7278 7644
rect 7214 7584 7278 7588
rect 7294 7644 7358 7648
rect 7294 7588 7298 7644
rect 7298 7588 7354 7644
rect 7354 7588 7358 7644
rect 7294 7584 7358 7588
rect 13157 7644 13221 7648
rect 13157 7588 13161 7644
rect 13161 7588 13217 7644
rect 13217 7588 13221 7644
rect 13157 7584 13221 7588
rect 13237 7644 13301 7648
rect 13237 7588 13241 7644
rect 13241 7588 13297 7644
rect 13297 7588 13301 7644
rect 13237 7584 13301 7588
rect 13317 7644 13381 7648
rect 13317 7588 13321 7644
rect 13321 7588 13377 7644
rect 13377 7588 13381 7644
rect 13317 7584 13381 7588
rect 13397 7644 13461 7648
rect 13397 7588 13401 7644
rect 13401 7588 13457 7644
rect 13457 7588 13461 7644
rect 13397 7584 13461 7588
rect 4003 7100 4067 7104
rect 4003 7044 4007 7100
rect 4007 7044 4063 7100
rect 4063 7044 4067 7100
rect 4003 7040 4067 7044
rect 4083 7100 4147 7104
rect 4083 7044 4087 7100
rect 4087 7044 4143 7100
rect 4143 7044 4147 7100
rect 4083 7040 4147 7044
rect 4163 7100 4227 7104
rect 4163 7044 4167 7100
rect 4167 7044 4223 7100
rect 4223 7044 4227 7100
rect 4163 7040 4227 7044
rect 4243 7100 4307 7104
rect 4243 7044 4247 7100
rect 4247 7044 4303 7100
rect 4303 7044 4307 7100
rect 4243 7040 4307 7044
rect 10106 7100 10170 7104
rect 10106 7044 10110 7100
rect 10110 7044 10166 7100
rect 10166 7044 10170 7100
rect 10106 7040 10170 7044
rect 10186 7100 10250 7104
rect 10186 7044 10190 7100
rect 10190 7044 10246 7100
rect 10246 7044 10250 7100
rect 10186 7040 10250 7044
rect 10266 7100 10330 7104
rect 10266 7044 10270 7100
rect 10270 7044 10326 7100
rect 10326 7044 10330 7100
rect 10266 7040 10330 7044
rect 10346 7100 10410 7104
rect 10346 7044 10350 7100
rect 10350 7044 10406 7100
rect 10406 7044 10410 7100
rect 10346 7040 10410 7044
rect 16208 7100 16272 7104
rect 16208 7044 16212 7100
rect 16212 7044 16268 7100
rect 16268 7044 16272 7100
rect 16208 7040 16272 7044
rect 16288 7100 16352 7104
rect 16288 7044 16292 7100
rect 16292 7044 16348 7100
rect 16348 7044 16352 7100
rect 16288 7040 16352 7044
rect 16368 7100 16432 7104
rect 16368 7044 16372 7100
rect 16372 7044 16428 7100
rect 16428 7044 16432 7100
rect 16368 7040 16432 7044
rect 16448 7100 16512 7104
rect 16448 7044 16452 7100
rect 16452 7044 16508 7100
rect 16508 7044 16512 7100
rect 16448 7040 16512 7044
rect 7054 6556 7118 6560
rect 7054 6500 7058 6556
rect 7058 6500 7114 6556
rect 7114 6500 7118 6556
rect 7054 6496 7118 6500
rect 7134 6556 7198 6560
rect 7134 6500 7138 6556
rect 7138 6500 7194 6556
rect 7194 6500 7198 6556
rect 7134 6496 7198 6500
rect 7214 6556 7278 6560
rect 7214 6500 7218 6556
rect 7218 6500 7274 6556
rect 7274 6500 7278 6556
rect 7214 6496 7278 6500
rect 7294 6556 7358 6560
rect 7294 6500 7298 6556
rect 7298 6500 7354 6556
rect 7354 6500 7358 6556
rect 7294 6496 7358 6500
rect 13157 6556 13221 6560
rect 13157 6500 13161 6556
rect 13161 6500 13217 6556
rect 13217 6500 13221 6556
rect 13157 6496 13221 6500
rect 13237 6556 13301 6560
rect 13237 6500 13241 6556
rect 13241 6500 13297 6556
rect 13297 6500 13301 6556
rect 13237 6496 13301 6500
rect 13317 6556 13381 6560
rect 13317 6500 13321 6556
rect 13321 6500 13377 6556
rect 13377 6500 13381 6556
rect 13317 6496 13381 6500
rect 13397 6556 13461 6560
rect 13397 6500 13401 6556
rect 13401 6500 13457 6556
rect 13457 6500 13461 6556
rect 13397 6496 13461 6500
rect 4003 6012 4067 6016
rect 4003 5956 4007 6012
rect 4007 5956 4063 6012
rect 4063 5956 4067 6012
rect 4003 5952 4067 5956
rect 4083 6012 4147 6016
rect 4083 5956 4087 6012
rect 4087 5956 4143 6012
rect 4143 5956 4147 6012
rect 4083 5952 4147 5956
rect 4163 6012 4227 6016
rect 4163 5956 4167 6012
rect 4167 5956 4223 6012
rect 4223 5956 4227 6012
rect 4163 5952 4227 5956
rect 4243 6012 4307 6016
rect 4243 5956 4247 6012
rect 4247 5956 4303 6012
rect 4303 5956 4307 6012
rect 4243 5952 4307 5956
rect 10106 6012 10170 6016
rect 10106 5956 10110 6012
rect 10110 5956 10166 6012
rect 10166 5956 10170 6012
rect 10106 5952 10170 5956
rect 10186 6012 10250 6016
rect 10186 5956 10190 6012
rect 10190 5956 10246 6012
rect 10246 5956 10250 6012
rect 10186 5952 10250 5956
rect 10266 6012 10330 6016
rect 10266 5956 10270 6012
rect 10270 5956 10326 6012
rect 10326 5956 10330 6012
rect 10266 5952 10330 5956
rect 10346 6012 10410 6016
rect 10346 5956 10350 6012
rect 10350 5956 10406 6012
rect 10406 5956 10410 6012
rect 10346 5952 10410 5956
rect 16208 6012 16272 6016
rect 16208 5956 16212 6012
rect 16212 5956 16268 6012
rect 16268 5956 16272 6012
rect 16208 5952 16272 5956
rect 16288 6012 16352 6016
rect 16288 5956 16292 6012
rect 16292 5956 16348 6012
rect 16348 5956 16352 6012
rect 16288 5952 16352 5956
rect 16368 6012 16432 6016
rect 16368 5956 16372 6012
rect 16372 5956 16428 6012
rect 16428 5956 16432 6012
rect 16368 5952 16432 5956
rect 16448 6012 16512 6016
rect 16448 5956 16452 6012
rect 16452 5956 16508 6012
rect 16508 5956 16512 6012
rect 16448 5952 16512 5956
rect 7054 5468 7118 5472
rect 7054 5412 7058 5468
rect 7058 5412 7114 5468
rect 7114 5412 7118 5468
rect 7054 5408 7118 5412
rect 7134 5468 7198 5472
rect 7134 5412 7138 5468
rect 7138 5412 7194 5468
rect 7194 5412 7198 5468
rect 7134 5408 7198 5412
rect 7214 5468 7278 5472
rect 7214 5412 7218 5468
rect 7218 5412 7274 5468
rect 7274 5412 7278 5468
rect 7214 5408 7278 5412
rect 7294 5468 7358 5472
rect 7294 5412 7298 5468
rect 7298 5412 7354 5468
rect 7354 5412 7358 5468
rect 7294 5408 7358 5412
rect 13157 5468 13221 5472
rect 13157 5412 13161 5468
rect 13161 5412 13217 5468
rect 13217 5412 13221 5468
rect 13157 5408 13221 5412
rect 13237 5468 13301 5472
rect 13237 5412 13241 5468
rect 13241 5412 13297 5468
rect 13297 5412 13301 5468
rect 13237 5408 13301 5412
rect 13317 5468 13381 5472
rect 13317 5412 13321 5468
rect 13321 5412 13377 5468
rect 13377 5412 13381 5468
rect 13317 5408 13381 5412
rect 13397 5468 13461 5472
rect 13397 5412 13401 5468
rect 13401 5412 13457 5468
rect 13457 5412 13461 5468
rect 13397 5408 13461 5412
rect 4003 4924 4067 4928
rect 4003 4868 4007 4924
rect 4007 4868 4063 4924
rect 4063 4868 4067 4924
rect 4003 4864 4067 4868
rect 4083 4924 4147 4928
rect 4083 4868 4087 4924
rect 4087 4868 4143 4924
rect 4143 4868 4147 4924
rect 4083 4864 4147 4868
rect 4163 4924 4227 4928
rect 4163 4868 4167 4924
rect 4167 4868 4223 4924
rect 4223 4868 4227 4924
rect 4163 4864 4227 4868
rect 4243 4924 4307 4928
rect 4243 4868 4247 4924
rect 4247 4868 4303 4924
rect 4303 4868 4307 4924
rect 4243 4864 4307 4868
rect 10106 4924 10170 4928
rect 10106 4868 10110 4924
rect 10110 4868 10166 4924
rect 10166 4868 10170 4924
rect 10106 4864 10170 4868
rect 10186 4924 10250 4928
rect 10186 4868 10190 4924
rect 10190 4868 10246 4924
rect 10246 4868 10250 4924
rect 10186 4864 10250 4868
rect 10266 4924 10330 4928
rect 10266 4868 10270 4924
rect 10270 4868 10326 4924
rect 10326 4868 10330 4924
rect 10266 4864 10330 4868
rect 10346 4924 10410 4928
rect 10346 4868 10350 4924
rect 10350 4868 10406 4924
rect 10406 4868 10410 4924
rect 10346 4864 10410 4868
rect 16208 4924 16272 4928
rect 16208 4868 16212 4924
rect 16212 4868 16268 4924
rect 16268 4868 16272 4924
rect 16208 4864 16272 4868
rect 16288 4924 16352 4928
rect 16288 4868 16292 4924
rect 16292 4868 16348 4924
rect 16348 4868 16352 4924
rect 16288 4864 16352 4868
rect 16368 4924 16432 4928
rect 16368 4868 16372 4924
rect 16372 4868 16428 4924
rect 16428 4868 16432 4924
rect 16368 4864 16432 4868
rect 16448 4924 16512 4928
rect 16448 4868 16452 4924
rect 16452 4868 16508 4924
rect 16508 4868 16512 4924
rect 16448 4864 16512 4868
rect 7054 4380 7118 4384
rect 7054 4324 7058 4380
rect 7058 4324 7114 4380
rect 7114 4324 7118 4380
rect 7054 4320 7118 4324
rect 7134 4380 7198 4384
rect 7134 4324 7138 4380
rect 7138 4324 7194 4380
rect 7194 4324 7198 4380
rect 7134 4320 7198 4324
rect 7214 4380 7278 4384
rect 7214 4324 7218 4380
rect 7218 4324 7274 4380
rect 7274 4324 7278 4380
rect 7214 4320 7278 4324
rect 7294 4380 7358 4384
rect 7294 4324 7298 4380
rect 7298 4324 7354 4380
rect 7354 4324 7358 4380
rect 7294 4320 7358 4324
rect 13157 4380 13221 4384
rect 13157 4324 13161 4380
rect 13161 4324 13217 4380
rect 13217 4324 13221 4380
rect 13157 4320 13221 4324
rect 13237 4380 13301 4384
rect 13237 4324 13241 4380
rect 13241 4324 13297 4380
rect 13297 4324 13301 4380
rect 13237 4320 13301 4324
rect 13317 4380 13381 4384
rect 13317 4324 13321 4380
rect 13321 4324 13377 4380
rect 13377 4324 13381 4380
rect 13317 4320 13381 4324
rect 13397 4380 13461 4384
rect 13397 4324 13401 4380
rect 13401 4324 13457 4380
rect 13457 4324 13461 4380
rect 13397 4320 13461 4324
rect 4003 3836 4067 3840
rect 4003 3780 4007 3836
rect 4007 3780 4063 3836
rect 4063 3780 4067 3836
rect 4003 3776 4067 3780
rect 4083 3836 4147 3840
rect 4083 3780 4087 3836
rect 4087 3780 4143 3836
rect 4143 3780 4147 3836
rect 4083 3776 4147 3780
rect 4163 3836 4227 3840
rect 4163 3780 4167 3836
rect 4167 3780 4223 3836
rect 4223 3780 4227 3836
rect 4163 3776 4227 3780
rect 4243 3836 4307 3840
rect 4243 3780 4247 3836
rect 4247 3780 4303 3836
rect 4303 3780 4307 3836
rect 4243 3776 4307 3780
rect 10106 3836 10170 3840
rect 10106 3780 10110 3836
rect 10110 3780 10166 3836
rect 10166 3780 10170 3836
rect 10106 3776 10170 3780
rect 10186 3836 10250 3840
rect 10186 3780 10190 3836
rect 10190 3780 10246 3836
rect 10246 3780 10250 3836
rect 10186 3776 10250 3780
rect 10266 3836 10330 3840
rect 10266 3780 10270 3836
rect 10270 3780 10326 3836
rect 10326 3780 10330 3836
rect 10266 3776 10330 3780
rect 10346 3836 10410 3840
rect 10346 3780 10350 3836
rect 10350 3780 10406 3836
rect 10406 3780 10410 3836
rect 10346 3776 10410 3780
rect 16208 3836 16272 3840
rect 16208 3780 16212 3836
rect 16212 3780 16268 3836
rect 16268 3780 16272 3836
rect 16208 3776 16272 3780
rect 16288 3836 16352 3840
rect 16288 3780 16292 3836
rect 16292 3780 16348 3836
rect 16348 3780 16352 3836
rect 16288 3776 16352 3780
rect 16368 3836 16432 3840
rect 16368 3780 16372 3836
rect 16372 3780 16428 3836
rect 16428 3780 16432 3836
rect 16368 3776 16432 3780
rect 16448 3836 16512 3840
rect 16448 3780 16452 3836
rect 16452 3780 16508 3836
rect 16508 3780 16512 3836
rect 16448 3776 16512 3780
rect 7054 3292 7118 3296
rect 7054 3236 7058 3292
rect 7058 3236 7114 3292
rect 7114 3236 7118 3292
rect 7054 3232 7118 3236
rect 7134 3292 7198 3296
rect 7134 3236 7138 3292
rect 7138 3236 7194 3292
rect 7194 3236 7198 3292
rect 7134 3232 7198 3236
rect 7214 3292 7278 3296
rect 7214 3236 7218 3292
rect 7218 3236 7274 3292
rect 7274 3236 7278 3292
rect 7214 3232 7278 3236
rect 7294 3292 7358 3296
rect 7294 3236 7298 3292
rect 7298 3236 7354 3292
rect 7354 3236 7358 3292
rect 7294 3232 7358 3236
rect 13157 3292 13221 3296
rect 13157 3236 13161 3292
rect 13161 3236 13217 3292
rect 13217 3236 13221 3292
rect 13157 3232 13221 3236
rect 13237 3292 13301 3296
rect 13237 3236 13241 3292
rect 13241 3236 13297 3292
rect 13297 3236 13301 3292
rect 13237 3232 13301 3236
rect 13317 3292 13381 3296
rect 13317 3236 13321 3292
rect 13321 3236 13377 3292
rect 13377 3236 13381 3292
rect 13317 3232 13381 3236
rect 13397 3292 13461 3296
rect 13397 3236 13401 3292
rect 13401 3236 13457 3292
rect 13457 3236 13461 3292
rect 13397 3232 13461 3236
rect 4003 2748 4067 2752
rect 4003 2692 4007 2748
rect 4007 2692 4063 2748
rect 4063 2692 4067 2748
rect 4003 2688 4067 2692
rect 4083 2748 4147 2752
rect 4083 2692 4087 2748
rect 4087 2692 4143 2748
rect 4143 2692 4147 2748
rect 4083 2688 4147 2692
rect 4163 2748 4227 2752
rect 4163 2692 4167 2748
rect 4167 2692 4223 2748
rect 4223 2692 4227 2748
rect 4163 2688 4227 2692
rect 4243 2748 4307 2752
rect 4243 2692 4247 2748
rect 4247 2692 4303 2748
rect 4303 2692 4307 2748
rect 4243 2688 4307 2692
rect 10106 2748 10170 2752
rect 10106 2692 10110 2748
rect 10110 2692 10166 2748
rect 10166 2692 10170 2748
rect 10106 2688 10170 2692
rect 10186 2748 10250 2752
rect 10186 2692 10190 2748
rect 10190 2692 10246 2748
rect 10246 2692 10250 2748
rect 10186 2688 10250 2692
rect 10266 2748 10330 2752
rect 10266 2692 10270 2748
rect 10270 2692 10326 2748
rect 10326 2692 10330 2748
rect 10266 2688 10330 2692
rect 10346 2748 10410 2752
rect 10346 2692 10350 2748
rect 10350 2692 10406 2748
rect 10406 2692 10410 2748
rect 10346 2688 10410 2692
rect 16208 2748 16272 2752
rect 16208 2692 16212 2748
rect 16212 2692 16268 2748
rect 16268 2692 16272 2748
rect 16208 2688 16272 2692
rect 16288 2748 16352 2752
rect 16288 2692 16292 2748
rect 16292 2692 16348 2748
rect 16348 2692 16352 2748
rect 16288 2688 16352 2692
rect 16368 2748 16432 2752
rect 16368 2692 16372 2748
rect 16372 2692 16428 2748
rect 16428 2692 16432 2748
rect 16368 2688 16432 2692
rect 16448 2748 16512 2752
rect 16448 2692 16452 2748
rect 16452 2692 16508 2748
rect 16508 2692 16512 2748
rect 16448 2688 16512 2692
rect 7054 2204 7118 2208
rect 7054 2148 7058 2204
rect 7058 2148 7114 2204
rect 7114 2148 7118 2204
rect 7054 2144 7118 2148
rect 7134 2204 7198 2208
rect 7134 2148 7138 2204
rect 7138 2148 7194 2204
rect 7194 2148 7198 2204
rect 7134 2144 7198 2148
rect 7214 2204 7278 2208
rect 7214 2148 7218 2204
rect 7218 2148 7274 2204
rect 7274 2148 7278 2204
rect 7214 2144 7278 2148
rect 7294 2204 7358 2208
rect 7294 2148 7298 2204
rect 7298 2148 7354 2204
rect 7354 2148 7358 2204
rect 7294 2144 7358 2148
rect 13157 2204 13221 2208
rect 13157 2148 13161 2204
rect 13161 2148 13217 2204
rect 13217 2148 13221 2204
rect 13157 2144 13221 2148
rect 13237 2204 13301 2208
rect 13237 2148 13241 2204
rect 13241 2148 13297 2204
rect 13297 2148 13301 2204
rect 13237 2144 13301 2148
rect 13317 2204 13381 2208
rect 13317 2148 13321 2204
rect 13321 2148 13377 2204
rect 13377 2148 13381 2204
rect 13317 2144 13381 2148
rect 13397 2204 13461 2208
rect 13397 2148 13401 2204
rect 13401 2148 13457 2204
rect 13457 2148 13461 2204
rect 13397 2144 13461 2148
<< metal4 >>
rect 3995 20160 4316 20176
rect 3995 20096 4003 20160
rect 4067 20096 4083 20160
rect 4147 20096 4163 20160
rect 4227 20096 4243 20160
rect 4307 20096 4316 20160
rect 3995 19072 4316 20096
rect 3995 19008 4003 19072
rect 4067 19008 4083 19072
rect 4147 19008 4163 19072
rect 4227 19008 4243 19072
rect 4307 19008 4316 19072
rect 3995 17984 4316 19008
rect 3995 17920 4003 17984
rect 4067 17920 4083 17984
rect 4147 17920 4163 17984
rect 4227 17920 4243 17984
rect 4307 17920 4316 17984
rect 3995 17206 4316 17920
rect 3995 16970 4037 17206
rect 4273 16970 4316 17206
rect 3995 16896 4316 16970
rect 3995 16832 4003 16896
rect 4067 16832 4083 16896
rect 4147 16832 4163 16896
rect 4227 16832 4243 16896
rect 4307 16832 4316 16896
rect 3995 15808 4316 16832
rect 3995 15744 4003 15808
rect 4067 15744 4083 15808
rect 4147 15744 4163 15808
rect 4227 15744 4243 15808
rect 4307 15744 4316 15808
rect 3995 14720 4316 15744
rect 3995 14656 4003 14720
rect 4067 14656 4083 14720
rect 4147 14656 4163 14720
rect 4227 14656 4243 14720
rect 4307 14656 4316 14720
rect 3995 13632 4316 14656
rect 3995 13568 4003 13632
rect 4067 13568 4083 13632
rect 4147 13568 4163 13632
rect 4227 13568 4243 13632
rect 4307 13568 4316 13632
rect 3995 12544 4316 13568
rect 3995 12480 4003 12544
rect 4067 12480 4083 12544
rect 4147 12480 4163 12544
rect 4227 12480 4243 12544
rect 4307 12480 4316 12544
rect 3995 11456 4316 12480
rect 3995 11392 4003 11456
rect 4067 11392 4083 11456
rect 4147 11392 4163 11456
rect 4227 11392 4243 11456
rect 4307 11392 4316 11456
rect 3995 11222 4316 11392
rect 3995 10986 4037 11222
rect 4273 10986 4316 11222
rect 3995 10368 4316 10986
rect 3995 10304 4003 10368
rect 4067 10304 4083 10368
rect 4147 10304 4163 10368
rect 4227 10304 4243 10368
rect 4307 10304 4316 10368
rect 3995 9280 4316 10304
rect 3995 9216 4003 9280
rect 4067 9216 4083 9280
rect 4147 9216 4163 9280
rect 4227 9216 4243 9280
rect 4307 9216 4316 9280
rect 3995 8192 4316 9216
rect 3995 8128 4003 8192
rect 4067 8128 4083 8192
rect 4147 8128 4163 8192
rect 4227 8128 4243 8192
rect 4307 8128 4316 8192
rect 3995 7104 4316 8128
rect 3995 7040 4003 7104
rect 4067 7040 4083 7104
rect 4147 7040 4163 7104
rect 4227 7040 4243 7104
rect 4307 7040 4316 7104
rect 3995 6016 4316 7040
rect 3995 5952 4003 6016
rect 4067 5952 4083 6016
rect 4147 5952 4163 6016
rect 4227 5952 4243 6016
rect 4307 5952 4316 6016
rect 3995 5238 4316 5952
rect 3995 5002 4037 5238
rect 4273 5002 4316 5238
rect 3995 4928 4316 5002
rect 3995 4864 4003 4928
rect 4067 4864 4083 4928
rect 4147 4864 4163 4928
rect 4227 4864 4243 4928
rect 4307 4864 4316 4928
rect 3995 3840 4316 4864
rect 3995 3776 4003 3840
rect 4067 3776 4083 3840
rect 4147 3776 4163 3840
rect 4227 3776 4243 3840
rect 4307 3776 4316 3840
rect 3995 2752 4316 3776
rect 3995 2688 4003 2752
rect 4067 2688 4083 2752
rect 4147 2688 4163 2752
rect 4227 2688 4243 2752
rect 4307 2688 4316 2752
rect 3995 2128 4316 2688
rect 7046 19616 7366 20176
rect 7046 19552 7054 19616
rect 7118 19552 7134 19616
rect 7198 19552 7214 19616
rect 7278 19552 7294 19616
rect 7358 19552 7366 19616
rect 7046 18528 7366 19552
rect 7046 18464 7054 18528
rect 7118 18464 7134 18528
rect 7198 18464 7214 18528
rect 7278 18464 7294 18528
rect 7358 18464 7366 18528
rect 7046 17440 7366 18464
rect 7046 17376 7054 17440
rect 7118 17376 7134 17440
rect 7198 17376 7214 17440
rect 7278 17376 7294 17440
rect 7358 17376 7366 17440
rect 7046 16352 7366 17376
rect 7046 16288 7054 16352
rect 7118 16288 7134 16352
rect 7198 16288 7214 16352
rect 7278 16288 7294 16352
rect 7358 16288 7366 16352
rect 7046 15264 7366 16288
rect 7046 15200 7054 15264
rect 7118 15200 7134 15264
rect 7198 15200 7214 15264
rect 7278 15200 7294 15264
rect 7358 15200 7366 15264
rect 7046 14214 7366 15200
rect 7046 14176 7088 14214
rect 7324 14176 7366 14214
rect 7046 14112 7054 14176
rect 7358 14112 7366 14176
rect 7046 13978 7088 14112
rect 7324 13978 7366 14112
rect 7046 13088 7366 13978
rect 7046 13024 7054 13088
rect 7118 13024 7134 13088
rect 7198 13024 7214 13088
rect 7278 13024 7294 13088
rect 7358 13024 7366 13088
rect 7046 12000 7366 13024
rect 7046 11936 7054 12000
rect 7118 11936 7134 12000
rect 7198 11936 7214 12000
rect 7278 11936 7294 12000
rect 7358 11936 7366 12000
rect 7046 10912 7366 11936
rect 7046 10848 7054 10912
rect 7118 10848 7134 10912
rect 7198 10848 7214 10912
rect 7278 10848 7294 10912
rect 7358 10848 7366 10912
rect 7046 9824 7366 10848
rect 7046 9760 7054 9824
rect 7118 9760 7134 9824
rect 7198 9760 7214 9824
rect 7278 9760 7294 9824
rect 7358 9760 7366 9824
rect 7046 8736 7366 9760
rect 7046 8672 7054 8736
rect 7118 8672 7134 8736
rect 7198 8672 7214 8736
rect 7278 8672 7294 8736
rect 7358 8672 7366 8736
rect 7046 8230 7366 8672
rect 7046 7994 7088 8230
rect 7324 7994 7366 8230
rect 7046 7648 7366 7994
rect 7046 7584 7054 7648
rect 7118 7584 7134 7648
rect 7198 7584 7214 7648
rect 7278 7584 7294 7648
rect 7358 7584 7366 7648
rect 7046 6560 7366 7584
rect 7046 6496 7054 6560
rect 7118 6496 7134 6560
rect 7198 6496 7214 6560
rect 7278 6496 7294 6560
rect 7358 6496 7366 6560
rect 7046 5472 7366 6496
rect 7046 5408 7054 5472
rect 7118 5408 7134 5472
rect 7198 5408 7214 5472
rect 7278 5408 7294 5472
rect 7358 5408 7366 5472
rect 7046 4384 7366 5408
rect 7046 4320 7054 4384
rect 7118 4320 7134 4384
rect 7198 4320 7214 4384
rect 7278 4320 7294 4384
rect 7358 4320 7366 4384
rect 7046 3296 7366 4320
rect 7046 3232 7054 3296
rect 7118 3232 7134 3296
rect 7198 3232 7214 3296
rect 7278 3232 7294 3296
rect 7358 3232 7366 3296
rect 7046 2208 7366 3232
rect 7046 2144 7054 2208
rect 7118 2144 7134 2208
rect 7198 2144 7214 2208
rect 7278 2144 7294 2208
rect 7358 2144 7366 2208
rect 7046 2128 7366 2144
rect 10098 20160 10418 20176
rect 10098 20096 10106 20160
rect 10170 20096 10186 20160
rect 10250 20096 10266 20160
rect 10330 20096 10346 20160
rect 10410 20096 10418 20160
rect 10098 19072 10418 20096
rect 10098 19008 10106 19072
rect 10170 19008 10186 19072
rect 10250 19008 10266 19072
rect 10330 19008 10346 19072
rect 10410 19008 10418 19072
rect 10098 17984 10418 19008
rect 10098 17920 10106 17984
rect 10170 17920 10186 17984
rect 10250 17920 10266 17984
rect 10330 17920 10346 17984
rect 10410 17920 10418 17984
rect 10098 17206 10418 17920
rect 10098 16970 10140 17206
rect 10376 16970 10418 17206
rect 10098 16896 10418 16970
rect 10098 16832 10106 16896
rect 10170 16832 10186 16896
rect 10250 16832 10266 16896
rect 10330 16832 10346 16896
rect 10410 16832 10418 16896
rect 10098 15808 10418 16832
rect 10098 15744 10106 15808
rect 10170 15744 10186 15808
rect 10250 15744 10266 15808
rect 10330 15744 10346 15808
rect 10410 15744 10418 15808
rect 10098 14720 10418 15744
rect 10098 14656 10106 14720
rect 10170 14656 10186 14720
rect 10250 14656 10266 14720
rect 10330 14656 10346 14720
rect 10410 14656 10418 14720
rect 10098 13632 10418 14656
rect 10098 13568 10106 13632
rect 10170 13568 10186 13632
rect 10250 13568 10266 13632
rect 10330 13568 10346 13632
rect 10410 13568 10418 13632
rect 10098 12544 10418 13568
rect 10098 12480 10106 12544
rect 10170 12480 10186 12544
rect 10250 12480 10266 12544
rect 10330 12480 10346 12544
rect 10410 12480 10418 12544
rect 10098 11456 10418 12480
rect 10098 11392 10106 11456
rect 10170 11392 10186 11456
rect 10250 11392 10266 11456
rect 10330 11392 10346 11456
rect 10410 11392 10418 11456
rect 10098 11222 10418 11392
rect 10098 10986 10140 11222
rect 10376 10986 10418 11222
rect 10098 10368 10418 10986
rect 10098 10304 10106 10368
rect 10170 10304 10186 10368
rect 10250 10304 10266 10368
rect 10330 10304 10346 10368
rect 10410 10304 10418 10368
rect 10098 9280 10418 10304
rect 10098 9216 10106 9280
rect 10170 9216 10186 9280
rect 10250 9216 10266 9280
rect 10330 9216 10346 9280
rect 10410 9216 10418 9280
rect 10098 8192 10418 9216
rect 10098 8128 10106 8192
rect 10170 8128 10186 8192
rect 10250 8128 10266 8192
rect 10330 8128 10346 8192
rect 10410 8128 10418 8192
rect 10098 7104 10418 8128
rect 10098 7040 10106 7104
rect 10170 7040 10186 7104
rect 10250 7040 10266 7104
rect 10330 7040 10346 7104
rect 10410 7040 10418 7104
rect 10098 6016 10418 7040
rect 10098 5952 10106 6016
rect 10170 5952 10186 6016
rect 10250 5952 10266 6016
rect 10330 5952 10346 6016
rect 10410 5952 10418 6016
rect 10098 5238 10418 5952
rect 10098 5002 10140 5238
rect 10376 5002 10418 5238
rect 10098 4928 10418 5002
rect 10098 4864 10106 4928
rect 10170 4864 10186 4928
rect 10250 4864 10266 4928
rect 10330 4864 10346 4928
rect 10410 4864 10418 4928
rect 10098 3840 10418 4864
rect 10098 3776 10106 3840
rect 10170 3776 10186 3840
rect 10250 3776 10266 3840
rect 10330 3776 10346 3840
rect 10410 3776 10418 3840
rect 10098 2752 10418 3776
rect 10098 2688 10106 2752
rect 10170 2688 10186 2752
rect 10250 2688 10266 2752
rect 10330 2688 10346 2752
rect 10410 2688 10418 2752
rect 10098 2128 10418 2688
rect 13149 19616 13469 20176
rect 13149 19552 13157 19616
rect 13221 19552 13237 19616
rect 13301 19552 13317 19616
rect 13381 19552 13397 19616
rect 13461 19552 13469 19616
rect 13149 18528 13469 19552
rect 13149 18464 13157 18528
rect 13221 18464 13237 18528
rect 13301 18464 13317 18528
rect 13381 18464 13397 18528
rect 13461 18464 13469 18528
rect 13149 17440 13469 18464
rect 13149 17376 13157 17440
rect 13221 17376 13237 17440
rect 13301 17376 13317 17440
rect 13381 17376 13397 17440
rect 13461 17376 13469 17440
rect 13149 16352 13469 17376
rect 13149 16288 13157 16352
rect 13221 16288 13237 16352
rect 13301 16288 13317 16352
rect 13381 16288 13397 16352
rect 13461 16288 13469 16352
rect 13149 15264 13469 16288
rect 13149 15200 13157 15264
rect 13221 15200 13237 15264
rect 13301 15200 13317 15264
rect 13381 15200 13397 15264
rect 13461 15200 13469 15264
rect 13149 14214 13469 15200
rect 13149 14176 13191 14214
rect 13427 14176 13469 14214
rect 13149 14112 13157 14176
rect 13461 14112 13469 14176
rect 13149 13978 13191 14112
rect 13427 13978 13469 14112
rect 13149 13088 13469 13978
rect 13149 13024 13157 13088
rect 13221 13024 13237 13088
rect 13301 13024 13317 13088
rect 13381 13024 13397 13088
rect 13461 13024 13469 13088
rect 13149 12000 13469 13024
rect 13149 11936 13157 12000
rect 13221 11936 13237 12000
rect 13301 11936 13317 12000
rect 13381 11936 13397 12000
rect 13461 11936 13469 12000
rect 13149 10912 13469 11936
rect 13149 10848 13157 10912
rect 13221 10848 13237 10912
rect 13301 10848 13317 10912
rect 13381 10848 13397 10912
rect 13461 10848 13469 10912
rect 13149 9824 13469 10848
rect 13149 9760 13157 9824
rect 13221 9760 13237 9824
rect 13301 9760 13317 9824
rect 13381 9760 13397 9824
rect 13461 9760 13469 9824
rect 13149 8736 13469 9760
rect 13149 8672 13157 8736
rect 13221 8672 13237 8736
rect 13301 8672 13317 8736
rect 13381 8672 13397 8736
rect 13461 8672 13469 8736
rect 13149 8230 13469 8672
rect 13149 7994 13191 8230
rect 13427 7994 13469 8230
rect 13149 7648 13469 7994
rect 13149 7584 13157 7648
rect 13221 7584 13237 7648
rect 13301 7584 13317 7648
rect 13381 7584 13397 7648
rect 13461 7584 13469 7648
rect 13149 6560 13469 7584
rect 13149 6496 13157 6560
rect 13221 6496 13237 6560
rect 13301 6496 13317 6560
rect 13381 6496 13397 6560
rect 13461 6496 13469 6560
rect 13149 5472 13469 6496
rect 13149 5408 13157 5472
rect 13221 5408 13237 5472
rect 13301 5408 13317 5472
rect 13381 5408 13397 5472
rect 13461 5408 13469 5472
rect 13149 4384 13469 5408
rect 13149 4320 13157 4384
rect 13221 4320 13237 4384
rect 13301 4320 13317 4384
rect 13381 4320 13397 4384
rect 13461 4320 13469 4384
rect 13149 3296 13469 4320
rect 13149 3232 13157 3296
rect 13221 3232 13237 3296
rect 13301 3232 13317 3296
rect 13381 3232 13397 3296
rect 13461 3232 13469 3296
rect 13149 2208 13469 3232
rect 13149 2144 13157 2208
rect 13221 2144 13237 2208
rect 13301 2144 13317 2208
rect 13381 2144 13397 2208
rect 13461 2144 13469 2208
rect 13149 2128 13469 2144
rect 16200 20160 16521 20176
rect 16200 20096 16208 20160
rect 16272 20096 16288 20160
rect 16352 20096 16368 20160
rect 16432 20096 16448 20160
rect 16512 20096 16521 20160
rect 16200 19072 16521 20096
rect 16200 19008 16208 19072
rect 16272 19008 16288 19072
rect 16352 19008 16368 19072
rect 16432 19008 16448 19072
rect 16512 19008 16521 19072
rect 16200 17984 16521 19008
rect 16200 17920 16208 17984
rect 16272 17920 16288 17984
rect 16352 17920 16368 17984
rect 16432 17920 16448 17984
rect 16512 17920 16521 17984
rect 16200 17206 16521 17920
rect 16200 16970 16242 17206
rect 16478 16970 16521 17206
rect 16200 16896 16521 16970
rect 16200 16832 16208 16896
rect 16272 16832 16288 16896
rect 16352 16832 16368 16896
rect 16432 16832 16448 16896
rect 16512 16832 16521 16896
rect 16200 15808 16521 16832
rect 16200 15744 16208 15808
rect 16272 15744 16288 15808
rect 16352 15744 16368 15808
rect 16432 15744 16448 15808
rect 16512 15744 16521 15808
rect 16200 14720 16521 15744
rect 16200 14656 16208 14720
rect 16272 14656 16288 14720
rect 16352 14656 16368 14720
rect 16432 14656 16448 14720
rect 16512 14656 16521 14720
rect 16200 13632 16521 14656
rect 16200 13568 16208 13632
rect 16272 13568 16288 13632
rect 16352 13568 16368 13632
rect 16432 13568 16448 13632
rect 16512 13568 16521 13632
rect 16200 12544 16521 13568
rect 16200 12480 16208 12544
rect 16272 12480 16288 12544
rect 16352 12480 16368 12544
rect 16432 12480 16448 12544
rect 16512 12480 16521 12544
rect 16200 11456 16521 12480
rect 16200 11392 16208 11456
rect 16272 11392 16288 11456
rect 16352 11392 16368 11456
rect 16432 11392 16448 11456
rect 16512 11392 16521 11456
rect 16200 11222 16521 11392
rect 16200 10986 16242 11222
rect 16478 10986 16521 11222
rect 16200 10368 16521 10986
rect 16200 10304 16208 10368
rect 16272 10304 16288 10368
rect 16352 10304 16368 10368
rect 16432 10304 16448 10368
rect 16512 10304 16521 10368
rect 16200 9280 16521 10304
rect 16200 9216 16208 9280
rect 16272 9216 16288 9280
rect 16352 9216 16368 9280
rect 16432 9216 16448 9280
rect 16512 9216 16521 9280
rect 16200 8192 16521 9216
rect 16200 8128 16208 8192
rect 16272 8128 16288 8192
rect 16352 8128 16368 8192
rect 16432 8128 16448 8192
rect 16512 8128 16521 8192
rect 16200 7104 16521 8128
rect 16200 7040 16208 7104
rect 16272 7040 16288 7104
rect 16352 7040 16368 7104
rect 16432 7040 16448 7104
rect 16512 7040 16521 7104
rect 16200 6016 16521 7040
rect 16200 5952 16208 6016
rect 16272 5952 16288 6016
rect 16352 5952 16368 6016
rect 16432 5952 16448 6016
rect 16512 5952 16521 6016
rect 16200 5238 16521 5952
rect 16200 5002 16242 5238
rect 16478 5002 16521 5238
rect 16200 4928 16521 5002
rect 16200 4864 16208 4928
rect 16272 4864 16288 4928
rect 16352 4864 16368 4928
rect 16432 4864 16448 4928
rect 16512 4864 16521 4928
rect 16200 3840 16521 4864
rect 16200 3776 16208 3840
rect 16272 3776 16288 3840
rect 16352 3776 16368 3840
rect 16432 3776 16448 3840
rect 16512 3776 16521 3840
rect 16200 2752 16521 3776
rect 16200 2688 16208 2752
rect 16272 2688 16288 2752
rect 16352 2688 16368 2752
rect 16432 2688 16448 2752
rect 16512 2688 16521 2752
rect 16200 2128 16521 2688
<< via4 >>
rect 4037 16970 4273 17206
rect 4037 10986 4273 11222
rect 4037 5002 4273 5238
rect 7088 14176 7324 14214
rect 7088 14112 7118 14176
rect 7118 14112 7134 14176
rect 7134 14112 7198 14176
rect 7198 14112 7214 14176
rect 7214 14112 7278 14176
rect 7278 14112 7294 14176
rect 7294 14112 7324 14176
rect 7088 13978 7324 14112
rect 7088 7994 7324 8230
rect 10140 16970 10376 17206
rect 10140 10986 10376 11222
rect 10140 5002 10376 5238
rect 13191 14176 13427 14214
rect 13191 14112 13221 14176
rect 13221 14112 13237 14176
rect 13237 14112 13301 14176
rect 13301 14112 13317 14176
rect 13317 14112 13381 14176
rect 13381 14112 13397 14176
rect 13397 14112 13427 14176
rect 13191 13978 13427 14112
rect 13191 7994 13427 8230
rect 16242 16970 16478 17206
rect 16242 10986 16478 11222
rect 16242 5002 16478 5238
<< metal5 >>
rect 1104 17206 19412 17248
rect 1104 16970 4037 17206
rect 4273 16970 10140 17206
rect 10376 16970 16242 17206
rect 16478 16970 19412 17206
rect 1104 16928 19412 16970
rect 1104 14214 19412 14256
rect 1104 13978 7088 14214
rect 7324 13978 13191 14214
rect 13427 13978 19412 14214
rect 1104 13936 19412 13978
rect 1104 11222 19412 11264
rect 1104 10986 4037 11222
rect 4273 10986 10140 11222
rect 10376 10986 16242 11222
rect 16478 10986 19412 11222
rect 1104 10944 19412 10986
rect 1104 8230 19412 8272
rect 1104 7994 7088 8230
rect 7324 7994 13191 8230
rect 13427 7994 19412 8230
rect 1104 7952 19412 7994
rect 1104 5238 19412 5280
rect 1104 5002 4037 5238
rect 4273 5002 10140 5238
rect 10376 5002 16242 5238
rect 16478 5002 19412 5238
rect 1104 4960 19412 5002
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 0
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_144
timestamp 0
transform 1 0 14352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 0
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 0
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18
timestamp 0
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 0
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 0
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_79
timestamp 0
transform 1 0 8372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 0
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 0
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 0
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_157
timestamp 0
transform 1 0 15548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 0
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 0
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 0
transform 1 0 18032 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 0
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_59
timestamp 0
transform 1 0 6532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_67
timestamp 0
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 0
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 0
transform 1 0 10764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_117
timestamp 0
transform 1 0 11868 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_131
timestamp 0
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 0
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 0
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_176
timestamp 0
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 0
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 0
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 0
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_24
timestamp 0
transform 1 0 3312 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 0
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_65
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 0
transform 1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_79
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_91
timestamp 0
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 0
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_121
timestamp 0
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_144
timestamp 0
transform 1 0 14352 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_148
timestamp 0
transform 1 0 14720 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 0
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_189
timestamp 0
transform 1 0 18492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_195
timestamp 0
transform 1 0 19044 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_16
timestamp 0
transform 1 0 2576 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_46
timestamp 0
transform 1 0 5336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_54
timestamp 0
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_64
timestamp 0
transform 1 0 6992 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 0
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 0
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 0
transform 1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_108
timestamp 0
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_120
timestamp 0
transform 1 0 12144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_127
timestamp 0
transform 1 0 12788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 0
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_146
timestamp 0
transform 1 0 14536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_157
timestamp 0
transform 1 0 15548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_169
timestamp 0
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_173
timestamp 0
transform 1 0 17020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 0
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_188
timestamp 0
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_11
timestamp 0
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 0
transform 1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 0
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_66
timestamp 0
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_74
timestamp 0
transform 1 0 7912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 0
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 0
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_116
timestamp 0
transform 1 0 11776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_127
timestamp 0
transform 1 0 12788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_134
timestamp 0
transform 1 0 13432 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 0
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_153
timestamp 0
transform 1 0 15180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 0
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_180
timestamp 0
transform 1 0 17664 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_189
timestamp 0
transform 1 0 18492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_195
timestamp 0
transform 1 0 19044 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 0
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_35
timestamp 0
transform 1 0 4324 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_48
timestamp 0
transform 1 0 5520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp 0
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_95
timestamp 0
transform 1 0 9844 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp 0
transform 1 0 10580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_129
timestamp 0
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 0
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_162
timestamp 0
transform 1 0 16008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 0
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 0
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_9
timestamp 0
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_21
timestamp 0
transform 1 0 3036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_29
timestamp 0
transform 1 0 3772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 0
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 0
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_60
timestamp 0
transform 1 0 6624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_68
timestamp 0
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_76
timestamp 0
transform 1 0 8096 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_88
timestamp 0
transform 1 0 9200 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_100
timestamp 0
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_133
timestamp 0
transform 1 0 13340 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 0
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 0
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_193
timestamp 0
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_49
timestamp 0
transform 1 0 5612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_61
timestamp 0
transform 1 0 6716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_67
timestamp 0
transform 1 0 7268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 0
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_95
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_107
timestamp 0
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_119
timestamp 0
transform 1 0 12052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 0
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 0
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_152
timestamp 0
transform 1 0 15088 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_176
timestamp 0
transform 1 0 17296 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_183
timestamp 0
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 0
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 0
transform 1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_26
timestamp 0
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_38
timestamp 0
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 0
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 0
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_88
timestamp 0
transform 1 0 9200 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_94
timestamp 0
transform 1 0 9752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 0
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 0
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_132
timestamp 0
transform 1 0 13248 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_142
timestamp 0
transform 1 0 14168 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 0
transform 1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 0
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 0
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_192
timestamp 0
transform 1 0 18768 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 0
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_37
timestamp 0
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_44
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 0
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 0
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 0
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 0
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 0
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 0
transform 1 0 12972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 0
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_161
timestamp 0
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_173
timestamp 0
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_181
timestamp 0
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 0
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 0
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 0
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 0
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 0
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_61
timestamp 0
transform 1 0 6716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_67
timestamp 0
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 0
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 0
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_92
timestamp 0
transform 1 0 9568 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_104
timestamp 0
transform 1 0 10672 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 0
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 0
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 0
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_152
timestamp 0
transform 1 0 15088 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 0
transform 1 0 15824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 0
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_176
timestamp 0
transform 1 0 17296 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 0
transform 1 0 17848 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_190
timestamp 0
transform 1 0 18584 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_35
timestamp 0
transform 1 0 4324 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 0
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_50
timestamp 0
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 0
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_72
timestamp 0
transform 1 0 7728 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 0
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 0
transform 1 0 10120 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_110
timestamp 0
transform 1 0 11224 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_120
timestamp 0
transform 1 0 12144 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 0
transform 1 0 12880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 0
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_145
timestamp 0
transform 1 0 14444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_149
timestamp 0
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 0
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_164
timestamp 0
transform 1 0 16192 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_179
timestamp 0
transform 1 0 17572 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 0
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_9
timestamp 0
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_21
timestamp 0
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_31
timestamp 0
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 0
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 0
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_77
timestamp 0
transform 1 0 8188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_85
timestamp 0
transform 1 0 8924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_95
timestamp 0
transform 1 0 9844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 0
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_121
timestamp 0
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_128
timestamp 0
transform 1 0 12880 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_154
timestamp 0
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 0
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 0
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_195
timestamp 0
transform 1 0 19044 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_10
timestamp 0
transform 1 0 2024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_16
timestamp 0
transform 1 0 2576 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 0
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_49
timestamp 0
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 0
transform 1 0 6348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 0
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 0
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 0
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 0
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 0
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 0
transform 1 0 14812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_160
timestamp 0
transform 1 0 15824 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 0
transform 1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 0
transform 1 0 17572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp 0
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 0
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_22
timestamp 0
transform 1 0 3128 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_34
timestamp 0
transform 1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_42
timestamp 0
transform 1 0 4968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_48
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 0
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 0
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_82
timestamp 0
transform 1 0 8648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_86
timestamp 0
transform 1 0 9016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_94
timestamp 0
transform 1 0 9752 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 0
transform 1 0 10304 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 0
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_118
timestamp 0
transform 1 0 11960 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 0
transform 1 0 14536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 0
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 0
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 0
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 0
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_37
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 0
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 0
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 0
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_92
timestamp 0
transform 1 0 9568 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 0
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_125
timestamp 0
transform 1 0 12604 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 0
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_146
timestamp 0
transform 1 0 14536 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 0
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 0
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 0
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_7
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_16
timestamp 0
transform 1 0 2576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_28
timestamp 0
transform 1 0 3680 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_36
timestamp 0
transform 1 0 4416 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_41
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 0
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_68
timestamp 0
transform 1 0 7360 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_76
timestamp 0
transform 1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 0
transform 1 0 10212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 0
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_120
timestamp 0
transform 1 0 12144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 0
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_132
timestamp 0
transform 1 0 13248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 0
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_155
timestamp 0
transform 1 0 15364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_172
timestamp 0
transform 1 0 16928 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_187
timestamp 0
transform 1 0 18308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_195
timestamp 0
transform 1 0 19044 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_49
timestamp 0
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_61
timestamp 0
transform 1 0 6716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 0
transform 1 0 10488 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_126
timestamp 0
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 0
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 0
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_156
timestamp 0
transform 1 0 15456 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_169
timestamp 0
transform 1 0 16652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_181
timestamp 0
transform 1 0 17756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 0
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 0
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_21
timestamp 0
transform 1 0 3036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 0
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_34
timestamp 0
transform 1 0 4232 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 0
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_64
timestamp 0
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 0
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_75
timestamp 0
transform 1 0 8004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_80
timestamp 0
transform 1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_87
timestamp 0
transform 1 0 9108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 0
transform 1 0 10120 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 0
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 0
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 0
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_138
timestamp 0
transform 1 0 13800 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_146
timestamp 0
transform 1 0 14536 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 0
transform 1 0 15088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 0
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_177
timestamp 0
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 0
transform 1 0 18032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 0
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_195
timestamp 0
transform 1 0 19044 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 0
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 0
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 0
transform 1 0 4048 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_44
timestamp 0
transform 1 0 5152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_48
timestamp 0
transform 1 0 5520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_56
timestamp 0
transform 1 0 6256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_64
timestamp 0
transform 1 0 6992 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_70
timestamp 0
transform 1 0 7544 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 0
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_98
timestamp 0
transform 1 0 10120 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_106
timestamp 0
transform 1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_116
timestamp 0
transform 1 0 11776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_128
timestamp 0
transform 1 0 12880 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 0
transform 1 0 14352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_152
timestamp 0
transform 1 0 15088 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_160
timestamp 0
transform 1 0 15824 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_168
timestamp 0
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 0
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 0
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 0
transform 1 0 4048 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp 0
transform 1 0 4416 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_41
timestamp 0
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 0
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_77
timestamp 0
transform 1 0 8188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_85
timestamp 0
transform 1 0 8924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 0
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 0
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 0
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_141
timestamp 0
transform 1 0 14076 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_154
timestamp 0
transform 1 0 15272 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 0
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 0
transform 1 0 16928 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 0
transform 1 0 18032 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 0
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 0
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 0
transform 1 0 5612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_57
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_72
timestamp 0
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_88
timestamp 0
transform 1 0 9200 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_96
timestamp 0
transform 1 0 9936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_106
timestamp 0
transform 1 0 10856 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 0
transform 1 0 11684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 0
transform 1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 0
transform 1 0 13156 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 0
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_161
timestamp 0
transform 1 0 15916 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_176
timestamp 0
transform 1 0 17296 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_182
timestamp 0
transform 1 0 17848 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 0
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_35
timestamp 0
transform 1 0 4324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 0
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 0
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_92
timestamp 0
transform 1 0 9568 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 0
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 0
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_121
timestamp 0
transform 1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_128
timestamp 0
transform 1 0 12880 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 0
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_147
timestamp 0
transform 1 0 14628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_158
timestamp 0
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 0
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_189
timestamp 0
transform 1 0 18492 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_195
timestamp 0
transform 1 0 19044 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 0
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 0
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 0
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_88
timestamp 0
transform 1 0 9200 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_96
timestamp 0
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 0
transform 1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_110
timestamp 0
transform 1 0 11224 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 0
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 0
transform 1 0 15088 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 0
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_174
timestamp 0
transform 1 0 17112 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 0
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 0
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 0
transform 1 0 2024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 0
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 0
transform 1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_37
timestamp 0
transform 1 0 4508 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_45
timestamp 0
transform 1 0 5244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_64
timestamp 0
transform 1 0 6992 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_92
timestamp 0
transform 1 0 9568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_103
timestamp 0
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_128
timestamp 0
transform 1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 0
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 0
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_156
timestamp 0
transform 1 0 15456 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_160
timestamp 0
transform 1 0 15824 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 0
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_176
timestamp 0
transform 1 0 17296 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 0
transform 1 0 17848 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_186
timestamp 0
transform 1 0 18216 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_194
timestamp 0
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 0
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_36
timestamp 0
transform 1 0 4416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_55
timestamp 0
transform 1 0 6164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 0
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 0
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_108
timestamp 0
transform 1 0 11040 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_116
timestamp 0
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_120
timestamp 0
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp 0
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_171
timestamp 0
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 0
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 0
transform 1 0 2852 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 0
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 0
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_77
timestamp 0
transform 1 0 8188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 0
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_90
timestamp 0
transform 1 0 9384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_99
timestamp 0
transform 1 0 10212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_133
timestamp 0
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 0
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_150
timestamp 0
transform 1 0 14904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 0
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_160
timestamp 0
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_173
timestamp 0
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 0
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_190
timestamp 0
transform 1 0 18584 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 0
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 0
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 0
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 0
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 0
transform 1 0 5244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_52
timestamp 0
transform 1 0 5888 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_59
timestamp 0
transform 1 0 6532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 0
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 0
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_105
timestamp 0
transform 1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_112
timestamp 0
transform 1 0 11408 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_125
timestamp 0
transform 1 0 12604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 0
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_146
timestamp 0
transform 1 0 14536 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 0
transform 1 0 15088 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 0
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 0
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_174
timestamp 0
transform 1 0 17112 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 0
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_24
timestamp 0
transform 1 0 3312 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 0
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_60
timestamp 0
transform 1 0 6624 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_71
timestamp 0
transform 1 0 7636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_83
timestamp 0
transform 1 0 8740 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_87
timestamp 0
transform 1 0 9108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 0
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 0
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_116
timestamp 0
transform 1 0 11776 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 0
transform 1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_130
timestamp 0
transform 1 0 13064 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_136
timestamp 0
transform 1 0 13616 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_140
timestamp 0
transform 1 0 13984 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_151
timestamp 0
transform 1 0 14996 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_159
timestamp 0
transform 1 0 15732 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 0
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_189
timestamp 0
transform 1 0 18492 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_195
timestamp 0
transform 1 0 19044 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 0
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 0
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_49
timestamp 0
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 0
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 0
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_95
timestamp 0
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_106
timestamp 0
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_113
timestamp 0
transform 1 0 11500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_124
timestamp 0
transform 1 0 12512 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 0
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 0
transform 1 0 15272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 0
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 0
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 0
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 0
transform 1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_27
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 0
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 0
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp 0
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_64
timestamp 0
transform 1 0 6992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_71
timestamp 0
transform 1 0 7636 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 0
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 0
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_135
timestamp 0
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 0
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 0
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_13
timestamp 0
transform 1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 0
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_37
timestamp 0
transform 1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_48
timestamp 0
transform 1 0 5520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_57
timestamp 0
transform 1 0 6348 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_69
timestamp 0
transform 1 0 7452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_95
timestamp 0
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_106
timestamp 0
transform 1 0 10856 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_123
timestamp 0
transform 1 0 12420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_131
timestamp 0
transform 1 0 13156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 0
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 0
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 0
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 0
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 0
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_190
timestamp 0
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 19412 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 19412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 19412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 19412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 19412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 19412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 19412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 19412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 19412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 19412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 6256 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 11408 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 16560 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _222_
timestamp 0
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _223_
timestamp 0
transform -1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _224_
timestamp 0
transform -1 0 2852 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _225_
timestamp 0
transform -1 0 3312 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _226_
timestamp 0
transform 1 0 1840 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _227_
timestamp 0
transform 1 0 14536 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _228_
timestamp 0
transform -1 0 12880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 0
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _230_
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _231_
timestamp 0
transform 1 0 14076 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 0
transform 1 0 13340 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _233_
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 0
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _235_
timestamp 0
transform -1 0 3312 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _236_
timestamp 0
transform 1 0 1840 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _237_
timestamp 0
transform 1 0 1932 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _238_
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _239_
timestamp 0
transform -1 0 2116 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _240_
timestamp 0
transform -1 0 5520 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _241_
timestamp 0
transform -1 0 5520 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _242_
timestamp 0
transform 1 0 3864 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _243_
timestamp 0
transform -1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _244_
timestamp 0
transform 1 0 4048 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _245_
timestamp 0
transform -1 0 4968 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _246_
timestamp 0
transform -1 0 4968 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _247_
timestamp 0
transform -1 0 3956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _248_
timestamp 0
transform -1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _249_
timestamp 0
transform 1 0 2668 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _250_
timestamp 0
transform -1 0 2852 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _251_
timestamp 0
transform -1 0 4048 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _252_
timestamp 0
transform 1 0 2300 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _253_
timestamp 0
transform 1 0 14720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _254_
timestamp 0
transform -1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _255_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _256_
timestamp 0
transform 1 0 2392 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _257_
timestamp 0
transform -1 0 5152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _258_
timestamp 0
transform 1 0 2392 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 0
transform 1 0 3404 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _260_
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _261_
timestamp 0
transform 1 0 4232 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _262_
timestamp 0
transform 1 0 2668 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _263_
timestamp 0
transform -1 0 3312 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _264_
timestamp 0
transform -1 0 4232 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _265_
timestamp 0
transform 1 0 2668 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 0
transform -1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _267_
timestamp 0
transform 1 0 2668 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _268_
timestamp 0
transform -1 0 7636 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _269_
timestamp 0
transform -1 0 8464 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _270_
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _271_
timestamp 0
transform -1 0 5520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _272_
timestamp 0
transform 1 0 4232 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _273_
timestamp 0
transform -1 0 8004 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _274_
timestamp 0
transform -1 0 7360 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _275_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _276_
timestamp 0
transform -1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _277_
timestamp 0
transform 1 0 5520 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _278_
timestamp 0
transform -1 0 7452 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _279_
timestamp 0
transform -1 0 7360 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _280_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _281_
timestamp 0
transform -1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _282_
timestamp 0
transform 1 0 7360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _283_
timestamp 0
transform 1 0 5612 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _284_
timestamp 0
transform -1 0 9660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _285_
timestamp 0
transform -1 0 7728 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _286_
timestamp 0
transform -1 0 7820 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _287_
timestamp 0
transform 1 0 6716 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 0
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _289_
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _290_
timestamp 0
transform -1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _291_
timestamp 0
transform -1 0 8096 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _292_
timestamp 0
transform 1 0 7268 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _293_
timestamp 0
transform -1 0 8464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _294_
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _295_
timestamp 0
transform -1 0 8280 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _296_
timestamp 0
transform -1 0 8372 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _297_
timestamp 0
transform 1 0 6624 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _298_
timestamp 0
transform -1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _299_
timestamp 0
transform 1 0 6348 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _300_
timestamp 0
transform -1 0 11040 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _301_
timestamp 0
transform -1 0 11132 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _302_
timestamp 0
transform 1 0 9200 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 0
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _304_
timestamp 0
transform 1 0 8096 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _305_
timestamp 0
transform -1 0 11040 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _306_
timestamp 0
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _307_
timestamp 0
transform 1 0 9200 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _308_
timestamp 0
transform -1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _309_
timestamp 0
transform -1 0 9568 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _310_
timestamp 0
transform 1 0 9108 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _311_
timestamp 0
transform -1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _312_
timestamp 0
transform -1 0 12972 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _313_
timestamp 0
transform -1 0 13800 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _314_
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _315_
timestamp 0
transform -1 0 10488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _316_
timestamp 0
transform 1 0 10396 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _317_
timestamp 0
transform 1 0 9200 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _318_
timestamp 0
transform 1 0 9660 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _319_
timestamp 0
transform 1 0 10212 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _320_
timestamp 0
transform -1 0 10396 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _321_
timestamp 0
transform 1 0 10212 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _322_
timestamp 0
transform 1 0 9384 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _323_
timestamp 0
transform 1 0 9752 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _324_
timestamp 0
transform 1 0 10396 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _325_
timestamp 0
transform -1 0 10488 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _326_
timestamp 0
transform -1 0 10580 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _327_
timestamp 0
transform -1 0 10856 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _328_
timestamp 0
transform 1 0 10580 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _329_
timestamp 0
transform 1 0 10212 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 0
transform -1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _331_
timestamp 0
transform 1 0 10120 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _332_
timestamp 0
transform -1 0 13156 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _333_
timestamp 0
transform -1 0 13432 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _334_
timestamp 0
transform 1 0 11960 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _335_
timestamp 0
transform -1 0 15272 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _336_
timestamp 0
transform 1 0 12880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _337_
timestamp 0
transform 1 0 11868 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 0
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _339_
timestamp 0
transform -1 0 15640 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _340_
timestamp 0
transform -1 0 15640 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _341_
timestamp 0
transform 1 0 13984 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _342_
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _343_
timestamp 0
transform -1 0 14720 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _344_
timestamp 0
transform -1 0 15272 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _345_
timestamp 0
transform -1 0 16100 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _346_
timestamp 0
transform 1 0 14352 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _347_
timestamp 0
transform -1 0 14536 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _348_
timestamp 0
transform 1 0 14260 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _349_
timestamp 0
transform -1 0 18584 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _350_
timestamp 0
transform -1 0 17572 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _351_
timestamp 0
transform -1 0 17112 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _352_
timestamp 0
transform -1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _353_
timestamp 0
transform 1 0 17940 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _354_
timestamp 0
transform -1 0 18584 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _355_
timestamp 0
transform -1 0 18584 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _356_
timestamp 0
transform 1 0 16652 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _357_
timestamp 0
transform -1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _358_
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _359_
timestamp 0
transform -1 0 18308 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _360_
timestamp 0
transform -1 0 18308 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _361_
timestamp 0
transform 1 0 16008 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _362_
timestamp 0
transform 1 0 17020 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _363_
timestamp 0
transform -1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _364_
timestamp 0
transform 1 0 15916 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _365_
timestamp 0
transform 1 0 14444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _366_
timestamp 0
transform 1 0 14904 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _367_
timestamp 0
transform -1 0 16100 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _368_
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _369_
timestamp 0
transform 1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _370_
timestamp 0
transform 1 0 15548 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _371_
timestamp 0
transform -1 0 18584 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _372_
timestamp 0
transform -1 0 18584 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _373_
timestamp 0
transform 1 0 16928 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _374_
timestamp 0
transform -1 0 16192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _375_
timestamp 0
transform -1 0 17296 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _376_
timestamp 0
transform 1 0 15364 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _377_
timestamp 0
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _378_
timestamp 0
transform 1 0 15640 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _379_
timestamp 0
transform -1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _380_
timestamp 0
transform 1 0 16652 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _381_
timestamp 0
transform -1 0 18308 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _382_
timestamp 0
transform -1 0 18032 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _383_
timestamp 0
transform 1 0 17112 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _384_
timestamp 0
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _385_
timestamp 0
transform -1 0 17664 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _386_
timestamp 0
transform 1 0 14352 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _387_
timestamp 0
transform 1 0 14720 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _388_
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _389_
timestamp 0
transform -1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _390_
timestamp 0
transform 1 0 14904 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _391_
timestamp 0
transform -1 0 13064 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _392_
timestamp 0
transform -1 0 13248 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _393_
timestamp 0
transform 1 0 12328 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _394_
timestamp 0
transform -1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _395_
timestamp 0
transform 1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _396_
timestamp 0
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _397_
timestamp 0
transform 1 0 12604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 0
transform -1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 0
transform -1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 0
transform 1 0 13156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 0
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _403_
timestamp 0
transform -1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _404_
timestamp 0
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 0
transform -1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 0
transform -1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 0
transform 1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 0
transform -1 0 5704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _410_
timestamp 0
transform -1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 0
transform -1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 0
transform 1 0 3956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 0
transform -1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 0
transform -1 0 4692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 0
transform -1 0 2300 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _416_
timestamp 0
transform -1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 0
transform -1 0 5244 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 0
transform 1 0 7360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 0
transform -1 0 5520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 0
transform 1 0 7452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 0
transform 1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _422_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 0
transform -1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 0
transform 1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 0
transform 1 0 6440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 0
transform -1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 0
transform 1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _428_
timestamp 0
transform -1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 0
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 0
transform -1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 0
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 0
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _434_
timestamp 0
transform -1 0 13432 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _435_
timestamp 0
transform -1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 0
transform -1 0 10120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 0
transform 1 0 11868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 0
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 0
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _441_
timestamp 0
transform -1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 0
transform 1 0 11408 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 0
transform -1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 0
transform -1 0 9200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 0
transform -1 0 9108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 0
transform 1 0 9108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _447_
timestamp 0
transform -1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 0
transform -1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 0
transform -1 0 13064 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 0
transform -1 0 13524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _453_
timestamp 0
transform 1 0 15640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 0
transform -1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 0
transform -1 0 15456 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 0
transform 1 0 17940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 0
transform 1 0 17480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 0
transform 1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _459_
timestamp 0
transform 1 0 14996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 0
transform 1 0 18400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 0
transform -1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 0
transform 1 0 17940 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 0
transform 1 0 17296 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _465_
timestamp 0
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 0
transform -1 0 15640 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 0
transform 1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 0
transform -1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 0
transform 1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 0
transform 1 0 18216 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 0
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 0
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 0
transform 1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _475_
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 0
transform -1 0 3220 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 0
transform -1 0 14536 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 0
transform -1 0 13616 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _479_
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _480_
timestamp 0
transform 1 0 1472 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _481_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 0
transform -1 0 5888 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 0
transform 1 0 3680 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _485_
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _486_
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _487_
timestamp 0
transform -1 0 3220 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 0
transform -1 0 5612 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 0
transform -1 0 3220 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 0
transform 1 0 5796 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 0
transform -1 0 5888 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 0
transform 1 0 5152 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 0
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _497_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _498_
timestamp 0
transform -1 0 8648 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _499_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 0
transform 1 0 6532 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 0
transform 1 0 6532 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _503_
timestamp 0
transform 1 0 9108 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp 0
transform -1 0 10764 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _505_
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 0
transform -1 0 12972 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 0
transform 1 0 10856 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _509_
timestamp 0
transform -1 0 10212 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _510_
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _511_
timestamp 0
transform 1 0 7728 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 0
transform 1 0 7728 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 0
transform -1 0 10212 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 0
transform -1 0 10764 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _515_
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 0
transform -1 0 13524 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _517_
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 0
transform 1 0 11500 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 0
transform 1 0 13892 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 0
transform 1 0 14444 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _521_
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _522_
timestamp 0
transform -1 0 18768 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _523_
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 0
transform 1 0 16928 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 0
transform 1 0 15640 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 0
transform 1 0 16928 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _527_
timestamp 0
transform 1 0 13432 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 0
transform 1 0 16928 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _529_
timestamp 0
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _530_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _531_
timestamp 0
transform 1 0 13892 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp 0
transform 1 0 16928 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _533_
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp 0
transform 1 0 16928 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _535_
timestamp 0
transform 1 0 12972 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp 0
transform 1 0 15456 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _537_
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _538_
timestamp 0
transform 1 0 12512 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 11960 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 0
transform -1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 0
transform 1 0 12512 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 0
transform -1 0 6348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 0
transform -1 0 6992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 0
transform -1 0 14076 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk
timestamp 0
transform -1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk
timestamp 0
transform 1 0 6532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk
timestamp 0
transform -1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk
timestamp 0
transform 1 0 6716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk
timestamp 0
transform -1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk
timestamp 0
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk
timestamp 0
transform -1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk
timestamp 0
transform 1 0 13248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 0
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 0
transform 1 0 6532 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 0
transform -1 0 8188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 0
transform 1 0 11500 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 11500 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 0
transform 1 0 12144 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 0
transform -1 0 12144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 0
transform -1 0 14168 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 0
transform -1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 0
transform -1 0 16284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 0
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 0
transform 1 0 16652 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 0
transform 1 0 16468 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 0
transform 1 0 17756 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 0
transform -1 0 16192 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 0
transform -1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 0
transform -1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 0
transform -1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 0
transform -1 0 18768 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 0
transform 1 0 2668 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 0
transform 1 0 4324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 0
transform -1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 0
transform 1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 0
transform -1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 0
transform -1 0 6532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 0
transform -1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 0
transform 1 0 13248 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
<< labels >>
rlabel metal5 s 1104 7952 19412 8272 4 VGND
port 1 nsew
rlabel metal5 s 1104 13936 19412 14256 4 VGND
port 1 nsew
rlabel metal4 s 7046 2128 7366 20176 4 VGND
port 1 nsew
rlabel metal4 s 13149 2128 13469 20176 4 VGND
port 1 nsew
rlabel metal5 s 1104 4960 19412 5280 4 VPWR
port 2 nsew
rlabel metal5 s 1104 10944 19412 11264 4 VPWR
port 2 nsew
rlabel metal5 s 1104 16928 19412 17248 4 VPWR
port 2 nsew
rlabel metal4 s 3996 2128 4316 20176 4 VPWR
port 2 nsew
rlabel metal4 s 10098 2128 10418 20176 4 VPWR
port 2 nsew
rlabel metal4 s 16201 2128 16521 20176 4 VPWR
port 2 nsew
rlabel metal3 s 19717 11296 20517 11416 4 clk
port 3 nsew
rlabel metal3 s 0 11296 800 11416 4 p
port 4 nsew
rlabel metal2 s 10230 0 10286 800 4 rst
port 5 nsew
rlabel metal2 s 294 21861 350 22661 4 x[0]
port 6 nsew
rlabel metal2 s 6458 21861 6514 22661 4 x[10]
port 7 nsew
rlabel metal2 s 7102 21861 7158 22661 4 x[11]
port 8 nsew
rlabel metal2 s 7746 21861 7802 22661 4 x[12]
port 9 nsew
rlabel metal2 s 8298 21861 8354 22661 4 x[13]
port 10 nsew
rlabel metal2 s 8942 21861 8998 22661 4 x[14]
port 11 nsew
rlabel metal2 s 9586 21861 9642 22661 4 x[15]
port 12 nsew
rlabel metal2 s 10230 21861 10286 22661 4 x[16]
port 13 nsew
rlabel metal2 s 10782 21861 10838 22661 4 x[17]
port 14 nsew
rlabel metal2 s 11426 21861 11482 22661 4 x[18]
port 15 nsew
rlabel metal2 s 12070 21861 12126 22661 4 x[19]
port 16 nsew
rlabel metal2 s 846 21861 902 22661 4 x[1]
port 17 nsew
rlabel metal2 s 12714 21861 12770 22661 4 x[20]
port 18 nsew
rlabel metal2 s 13266 21861 13322 22661 4 x[21]
port 19 nsew
rlabel metal2 s 13910 21861 13966 22661 4 x[22]
port 20 nsew
rlabel metal2 s 14554 21861 14610 22661 4 x[23]
port 21 nsew
rlabel metal2 s 15198 21861 15254 22661 4 x[24]
port 22 nsew
rlabel metal2 s 15750 21861 15806 22661 4 x[25]
port 23 nsew
rlabel metal2 s 16394 21861 16450 22661 4 x[26]
port 24 nsew
rlabel metal2 s 17038 21861 17094 22661 4 x[27]
port 25 nsew
rlabel metal2 s 17682 21861 17738 22661 4 x[28]
port 26 nsew
rlabel metal2 s 18234 21861 18290 22661 4 x[29]
port 27 nsew
rlabel metal2 s 1490 21861 1546 22661 4 x[2]
port 28 nsew
rlabel metal2 s 18878 21861 18934 22661 4 x[30]
port 29 nsew
rlabel metal2 s 19522 21861 19578 22661 4 x[31]
port 30 nsew
rlabel metal2 s 2134 21861 2190 22661 4 x[3]
port 31 nsew
rlabel metal2 s 2778 21861 2834 22661 4 x[4]
port 32 nsew
rlabel metal2 s 3330 21861 3386 22661 4 x[5]
port 33 nsew
rlabel metal2 s 3974 21861 4030 22661 4 x[6]
port 34 nsew
rlabel metal2 s 4618 21861 4674 22661 4 x[7]
port 35 nsew
rlabel metal2 s 5262 21861 5318 22661 4 x[8]
port 36 nsew
rlabel metal2 s 5814 21861 5870 22661 4 x[9]
port 37 nsew
rlabel metal2 s 20166 21861 20222 22661 4 y
port 38 nsew
<< properties >>
string FIXED_BBOX 0 0 20517 22661
<< end >>
