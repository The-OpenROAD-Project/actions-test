* NGSPICE file created from spm.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

.subckt spm VGND VPWR clk p rst x[0] x[10] x[11] x[12] x[13] x[14] x[15] x[16] x[17]
+ x[18] x[19] x[1] x[20] x[21] x[22] x[23] x[24] x[25] x[26] x[27] x[28] x[29] x[2]
+ x[30] x[31] x[3] x[4] x[5] x[6] x[7] x[8] x[9] y
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_363_ _384_/A _363_/B VGND VGND VPWR VPWR _364_/A sky130_fd_sc_hd__nand2_1
X_501_ _505_/CLK _501_/D _430_/Y VGND VGND VPWR VPWR _501_/Q sky130_fd_sc_hd__dfrtp_1
X_432_ _433_/A VGND VGND VPWR VPWR _432_/Y sky130_fd_sc_hd__inv_2
X_294_ _294_/A _294_/B VGND VGND VPWR VPWR _500_/D sky130_fd_sc_hd__xnor2_1
X_346_ _338_/X _347_/B _348_/B _345_/X VGND VGND VPWR VPWR _519_/D sky130_fd_sc_hd__a31o_1
X_415_ _415_/A VGND VGND VPWR VPWR _415_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_277_ _277_/A _277_/B VGND VGND VPWR VPWR _494_/D sky130_fd_sc_hd__xnor2_1
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_329_ _311_/X _330_/B _331_/B _328_/X VGND VGND VPWR VPWR _513_/D sky130_fd_sc_hd__a31o_1
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR _505_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_362_ _362_/A VGND VGND VPWR VPWR _384_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ _303_/A _293_/B VGND VGND VPWR VPWR _294_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_431_ _433_/A VGND VGND VPWR VPWR _431_/Y sky130_fd_sc_hd__inv_2
X_500_ _505_/CLK _500_/D _429_/Y VGND VGND VPWR VPWR _500_/Q sky130_fd_sc_hd__dfrtp_1
X_345_ _519_/Q _522_/Q VGND VGND VPWR VPWR _345_/X sky130_fd_sc_hd__and2_1
X_276_ _276_/A _276_/B VGND VGND VPWR VPWR _277_/A sky130_fd_sc_hd__nand2_1
X_414_ _415_/A VGND VGND VPWR VPWR _414_/Y sky130_fd_sc_hd__inv_2
X_328_ _513_/Q _516_/Q VGND VGND VPWR VPWR _328_/X sky130_fd_sc_hd__and2_1
X_259_ _487_/Q _490_/Q VGND VGND VPWR VPWR _259_/X sky130_fd_sc_hd__and2_1
XFILLER_2_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR _497_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_361_ _338_/X _363_/B _364_/B _360_/X VGND VGND VPWR VPWR _525_/D sky130_fd_sc_hd__a31o_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_430_ _433_/A VGND VGND VPWR VPWR _430_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_292_ _284_/X _293_/B _294_/B _291_/X VGND VGND VPWR VPWR _499_/D sky130_fd_sc_hd__a31o_1
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_344_ _519_/Q _522_/Q VGND VGND VPWR VPWR _348_/B sky130_fd_sc_hd__xor2_1
X_275_ _257_/X _276_/B _277_/B _274_/X VGND VGND VPWR VPWR _493_/D sky130_fd_sc_hd__a31o_1
X_413_ _415_/A VGND VGND VPWR VPWR _413_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_327_ _513_/Q _516_/Q VGND VGND VPWR VPWR _331_/B sky130_fd_sc_hd__xor2_1
X_258_ _487_/Q _490_/Q VGND VGND VPWR VPWR _262_/B sky130_fd_sc_hd__xor2_1
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_360_ _525_/Q _528_/Q VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__and2_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_291_ _499_/Q _502_/Q VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__and2_1
X_489_ _512_/CLK _489_/D _415_/Y VGND VGND VPWR VPWR _489_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ _343_/A _343_/B VGND VGND VPWR VPWR _518_/D sky130_fd_sc_hd__xnor2_1
X_274_ _493_/Q _496_/Q VGND VGND VPWR VPWR _274_/X sky130_fd_sc_hd__and2_1
X_412_ _415_/A VGND VGND VPWR VPWR _412_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_326_ _326_/A _326_/B VGND VGND VPWR VPWR _512_/D sky130_fd_sc_hd__xnor2_1
X_257_ _394_/A VGND VGND VPWR VPWR _257_/X sky130_fd_sc_hd__clkbuf_2
X_309_ _330_/A _309_/B VGND VGND VPWR VPWR _310_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_488_ _493_/CLK _488_/D _414_/Y VGND VGND VPWR VPWR _488_/Q sky130_fd_sc_hd__dfrtp_1
X_290_ _499_/Q _502_/Q VGND VGND VPWR VPWR _294_/B sky130_fd_sc_hd__xor2_1
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_273_ _493_/Q _496_/Q VGND VGND VPWR VPWR _277_/B sky130_fd_sc_hd__xor2_1
X_342_ _357_/A _342_/B VGND VGND VPWR VPWR _343_/A sky130_fd_sc_hd__nand2_1
X_411_ _415_/A VGND VGND VPWR VPWR _411_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ _330_/A _325_/B VGND VGND VPWR VPWR _326_/A sky130_fd_sc_hd__nand2_1
X_256_ _256_/A _256_/B VGND VGND VPWR VPWR _486_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_308_ _362_/A VGND VGND VPWR VPWR _330_/A sky130_fd_sc_hd__clkbuf_2
X_239_ _239_/A _239_/B VGND VGND VPWR VPWR _480_/D sky130_fd_sc_hd__xnor2_1
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput35 _476_/Q VGND VGND VPWR VPWR p sky130_fd_sc_hd__buf_2
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_487_ _493_/CLK _487_/D _413_/Y VGND VGND VPWR VPWR _487_/Q sky130_fd_sc_hd__dfrtp_1
X_272_ _272_/A _272_/B VGND VGND VPWR VPWR _492_/D sky130_fd_sc_hd__xnor2_1
X_341_ _338_/X _342_/B _343_/B _340_/X VGND VGND VPWR VPWR _517_/D sky130_fd_sc_hd__a31o_1
X_410_ _428_/A VGND VGND VPWR VPWR _415_/A sky130_fd_sc_hd__buf_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_324_ _311_/X _325_/B _326_/B _323_/X VGND VGND VPWR VPWR _511_/D sky130_fd_sc_hd__a31o_1
X_255_ _276_/A _255_/B VGND VGND VPWR VPWR _256_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_307_ _284_/X _309_/B _310_/B _306_/X VGND VGND VPWR VPWR _505_/D sky130_fd_sc_hd__a31o_1
X_238_ _248_/A _238_/B VGND VGND VPWR VPWR _239_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_486_ _493_/CLK _486_/D _412_/Y VGND VGND VPWR VPWR _486_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_271_ _276_/A _271_/B VGND VGND VPWR VPWR _272_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_340_ _517_/Q _520_/Q VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__and2_1
X_538_ _538_/CLK _538_/D _474_/Y VGND VGND VPWR VPWR _538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_469_ _470_/A VGND VGND VPWR VPWR _469_/Y sky130_fd_sc_hd__inv_2
X_323_ _511_/Q _514_/Q VGND VGND VPWR VPWR _323_/X sky130_fd_sc_hd__and2_1
X_254_ _362_/A VGND VGND VPWR VPWR _276_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_306_ _505_/Q _508_/Q VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__and2_1
X_237_ _223_/X _238_/B _239_/B _236_/X VGND VGND VPWR VPWR _479_/D sky130_fd_sc_hd__a31o_1
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_485_ _493_/CLK _485_/D _411_/Y VGND VGND VPWR VPWR _485_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_270_ _257_/X _271_/B _272_/B _269_/X VGND VGND VPWR VPWR _491_/D sky130_fd_sc_hd__a31o_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_399_ _402_/A VGND VGND VPWR VPWR _399_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_537_ _538_/CLK _537_/D _473_/Y VGND VGND VPWR VPWR _537_/Q sky130_fd_sc_hd__dfrtp_1
X_468_ _470_/A VGND VGND VPWR VPWR _468_/Y sky130_fd_sc_hd__inv_2
X_322_ _511_/Q _514_/Q VGND VGND VPWR VPWR _326_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_253_ _253_/A VGND VGND VPWR VPWR _362_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ _505_/Q _508_/Q VGND VGND VPWR VPWR _310_/B sky130_fd_sc_hd__xor2_1
X_236_ _479_/Q _482_/Q VGND VGND VPWR VPWR _236_/X sky130_fd_sc_hd__and2_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_484_ _497_/CLK _484_/D _409_/Y VGND VGND VPWR VPWR _484_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_536_ _536_/CLK _536_/D _472_/Y VGND VGND VPWR VPWR _536_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_467_ _470_/A VGND VGND VPWR VPWR _467_/Y sky130_fd_sc_hd__inv_2
X_398_ _402_/A VGND VGND VPWR VPWR _398_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_321_ _321_/A _321_/B VGND VGND VPWR VPWR _510_/D sky130_fd_sc_hd__xnor2_1
X_252_ _223_/X _255_/B _256_/B _251_/X VGND VGND VPWR VPWR _485_/D sky130_fd_sc_hd__a31o_1
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_519_ _526_/CLK _519_/D _452_/Y VGND VGND VPWR VPWR _519_/Q sky130_fd_sc_hd__dfrtp_1
X_235_ _479_/Q _482_/Q VGND VGND VPWR VPWR _239_/B sky130_fd_sc_hd__xor2_1
X_304_ _304_/A _304_/B VGND VGND VPWR VPWR _504_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_483_ _497_/CLK _483_/D _408_/Y VGND VGND VPWR VPWR _483_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_397_ _474_/A VGND VGND VPWR VPWR _402_/A sky130_fd_sc_hd__clkbuf_4
X_535_ _538_/CLK _535_/D _471_/Y VGND VGND VPWR VPWR _535_/Q sky130_fd_sc_hd__dfrtp_1
X_466_ _470_/A VGND VGND VPWR VPWR _466_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_320_ _330_/A _320_/B VGND VGND VPWR VPWR _321_/A sky130_fd_sc_hd__nand2_1
X_251_ _485_/Q _488_/Q VGND VGND VPWR VPWR _251_/X sky130_fd_sc_hd__and2_1
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_449_ _452_/A VGND VGND VPWR VPWR _449_/Y sky130_fd_sc_hd__inv_2
X_518_ _518_/CLK _518_/D _451_/Y VGND VGND VPWR VPWR _518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_234_ _234_/A VGND VGND VPWR VPWR _478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_303_ _303_/A _303_/B VGND VGND VPWR VPWR _304_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_482_ _505_/CLK _482_/D _407_/Y VGND VGND VPWR VPWR _482_/Q sky130_fd_sc_hd__dfrtp_1
X_396_ _465_/A VGND VGND VPWR VPWR _474_/A sky130_fd_sc_hd__clkbuf_2
X_534_ _536_/CLK _534_/D _470_/Y VGND VGND VPWR VPWR _534_/Q sky130_fd_sc_hd__dfrtp_1
X_465_ _465_/A VGND VGND VPWR VPWR _470_/A sky130_fd_sc_hd__buf_2
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_250_ _485_/Q _488_/Q VGND VGND VPWR VPWR _256_/B sky130_fd_sc_hd__xor2_1
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_448_ _452_/A VGND VGND VPWR VPWR _448_/Y sky130_fd_sc_hd__inv_2
X_517_ _526_/CLK _517_/D _450_/Y VGND VGND VPWR VPWR _517_/Q sky130_fd_sc_hd__dfrtp_1
X_379_ _384_/A _379_/B VGND VGND VPWR VPWR _380_/A sky130_fd_sc_hd__nand2_1
X_233_ _477_/D _233_/B VGND VGND VPWR VPWR _234_/A sky130_fd_sc_hd__and2_1
X_302_ _284_/X _303_/B _304_/B _301_/X VGND VGND VPWR VPWR _503_/D sky130_fd_sc_hd__a31o_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_481_ _497_/CLK _481_/D _406_/Y VGND VGND VPWR VPWR _481_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_464_ _464_/A VGND VGND VPWR VPWR _464_/Y sky130_fd_sc_hd__inv_2
X_533_ _536_/CLK _533_/D _469_/Y VGND VGND VPWR VPWR _533_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_395_ _395_/A _395_/B VGND VGND VPWR VPWR _538_/D sky130_fd_sc_hd__xnor2_1
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_516_ _526_/CLK _516_/D _449_/Y VGND VGND VPWR VPWR _516_/Q sky130_fd_sc_hd__dfrtp_1
X_447_ _459_/A VGND VGND VPWR VPWR _452_/A sky130_fd_sc_hd__buf_2
X_378_ _365_/X _379_/B _380_/B _377_/X VGND VGND VPWR VPWR _531_/D sky130_fd_sc_hd__a31o_1
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_232_ _365_/A _232_/B _477_/Q VGND VGND VPWR VPWR _233_/B sky130_fd_sc_hd__nand3_1
X_301_ _503_/Q _506_/Q VGND VGND VPWR VPWR _301_/X sky130_fd_sc_hd__and2_1
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_480_ _497_/CLK _480_/D _405_/Y VGND VGND VPWR VPWR _480_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_463_ _464_/A VGND VGND VPWR VPWR _463_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_394_ _394_/A _394_/B VGND VGND VPWR VPWR _395_/A sky130_fd_sc_hd__nand2_1
X_532_ _536_/CLK _532_/D _468_/Y VGND VGND VPWR VPWR _532_/Q sky130_fd_sc_hd__dfrtp_1
X_515_ _518_/CLK _515_/D _448_/Y VGND VGND VPWR VPWR _515_/Q sky130_fd_sc_hd__dfrtp_1
X_446_ _446_/A VGND VGND VPWR VPWR _446_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_377_ _531_/Q _534_/Q VGND VGND VPWR VPWR _377_/X sky130_fd_sc_hd__and2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_231_ _253_/A _232_/B _477_/Q VGND VGND VPWR VPWR _477_/D sky130_fd_sc_hd__a21o_1
X_300_ _503_/Q _506_/Q VGND VGND VPWR VPWR _304_/B sky130_fd_sc_hd__xor2_1
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_429_ _433_/A VGND VGND VPWR VPWR _429_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 rst VGND VGND VPWR VPWR _465_/A sky130_fd_sc_hd__clkbuf_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_393_ _248_/A _394_/B _395_/B _392_/X VGND VGND VPWR VPWR _537_/D sky130_fd_sc_hd__a31o_1
X_531_ _538_/CLK _531_/D _467_/Y VGND VGND VPWR VPWR _531_/Q sky130_fd_sc_hd__dfrtp_1
X_462_ _464_/A VGND VGND VPWR VPWR _462_/Y sky130_fd_sc_hd__inv_2
X_514_ _518_/CLK _514_/D _446_/Y VGND VGND VPWR VPWR _514_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_445_ _446_/A VGND VGND VPWR VPWR _445_/Y sky130_fd_sc_hd__inv_2
X_376_ _531_/Q _534_/Q VGND VGND VPWR VPWR _380_/B sky130_fd_sc_hd__xor2_1
X_230_ _230_/A _230_/B VGND VGND VPWR VPWR _476_/D sky130_fd_sc_hd__xnor2_1
X_359_ _525_/Q _528_/Q VGND VGND VPWR VPWR _364_/B sky130_fd_sc_hd__xor2_1
X_428_ _428_/A VGND VGND VPWR VPWR _433_/A sky130_fd_sc_hd__buf_2
Xinput2 x[0] VGND VGND VPWR VPWR _229_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_461_ _464_/A VGND VGND VPWR VPWR _461_/Y sky130_fd_sc_hd__inv_2
X_392_ _537_/Q _478_/Q VGND VGND VPWR VPWR _392_/X sky130_fd_sc_hd__and2_1
X_530_ _536_/CLK _530_/D _466_/Y VGND VGND VPWR VPWR _530_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_513_ _518_/CLK _513_/D _445_/Y VGND VGND VPWR VPWR _513_/Q sky130_fd_sc_hd__dfrtp_1
X_444_ _446_/A VGND VGND VPWR VPWR _444_/Y sky130_fd_sc_hd__inv_2
X_375_ _375_/A _375_/B VGND VGND VPWR VPWR _530_/D sky130_fd_sc_hd__xnor2_1
X_358_ _358_/A _358_/B VGND VGND VPWR VPWR _524_/D sky130_fd_sc_hd__xnor2_1
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_427_ _427_/A VGND VGND VPWR VPWR _427_/Y sky130_fd_sc_hd__inv_2
Xinput3 x[10] VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_289_ _289_/A _289_/B VGND VGND VPWR VPWR _498_/D sky130_fd_sc_hd__xnor2_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_460_ _464_/A VGND VGND VPWR VPWR _460_/Y sky130_fd_sc_hd__inv_2
X_391_ _537_/Q _478_/Q VGND VGND VPWR VPWR _395_/B sky130_fd_sc_hd__xor2_1
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_443_ _446_/A VGND VGND VPWR VPWR _443_/Y sky130_fd_sc_hd__inv_2
X_512_ _512_/CLK _512_/D _444_/Y VGND VGND VPWR VPWR _512_/Q sky130_fd_sc_hd__dfrtp_1
X_374_ _384_/A _374_/B VGND VGND VPWR VPWR _375_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 x[11] VGND VGND VPWR VPWR _293_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_357_ _357_/A _357_/B VGND VGND VPWR VPWR _358_/A sky130_fd_sc_hd__nand2_1
X_426_ _427_/A VGND VGND VPWR VPWR _426_/Y sky130_fd_sc_hd__inv_2
X_288_ _303_/A _288_/B VGND VGND VPWR VPWR _289_/A sky130_fd_sc_hd__nand2_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_409_ _409_/A VGND VGND VPWR VPWR _409_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_390_ _390_/A _390_/B VGND VGND VPWR VPWR _536_/D sky130_fd_sc_hd__xnor2_1
XFILLER_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_511_ _512_/CLK _511_/D _443_/Y VGND VGND VPWR VPWR _511_/Q sky130_fd_sc_hd__dfrtp_1
X_442_ _446_/A VGND VGND VPWR VPWR _442_/Y sky130_fd_sc_hd__inv_2
X_373_ _365_/X _374_/B _375_/B _372_/X VGND VGND VPWR VPWR _529_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 x[12] VGND VGND VPWR VPWR _298_/B sky130_fd_sc_hd__clkbuf_2
X_356_ _338_/X _357_/B _358_/B _355_/X VGND VGND VPWR VPWR _523_/D sky130_fd_sc_hd__a31o_1
X_287_ _284_/X _288_/B _289_/B _286_/X VGND VGND VPWR VPWR _497_/D sky130_fd_sc_hd__a31o_1
X_425_ _427_/A VGND VGND VPWR VPWR _425_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_408_ _409_/A VGND VGND VPWR VPWR _408_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_339_ _517_/Q _520_/Q VGND VGND VPWR VPWR _343_/B sky130_fd_sc_hd__xor2_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput30 x[6] VGND VGND VPWR VPWR _266_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_441_ _459_/A VGND VGND VPWR VPWR _446_/A sky130_fd_sc_hd__buf_2
X_510_ _518_/CLK _510_/D _442_/Y VGND VGND VPWR VPWR _510_/Q sky130_fd_sc_hd__dfrtp_1
X_372_ _529_/Q _532_/Q VGND VGND VPWR VPWR _372_/X sky130_fd_sc_hd__and2_1
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_355_ _523_/Q _526_/Q VGND VGND VPWR VPWR _355_/X sky130_fd_sc_hd__and2_1
X_424_ _427_/A VGND VGND VPWR VPWR _424_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_286_ _497_/Q _500_/Q VGND VGND VPWR VPWR _286_/X sky130_fd_sc_hd__and2_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput6 x[13] VGND VGND VPWR VPWR _303_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_269_ _491_/Q _494_/Q VGND VGND VPWR VPWR _269_/X sky130_fd_sc_hd__and2_1
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_338_ _365_/A VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__clkbuf_2
X_407_ _409_/A VGND VGND VPWR VPWR _407_/Y sky130_fd_sc_hd__inv_2
Xinput20 x[26] VGND VGND VPWR VPWR _374_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput31 x[7] VGND VGND VPWR VPWR _271_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_440_ _440_/A VGND VGND VPWR VPWR _440_/Y sky130_fd_sc_hd__inv_2
X_371_ _529_/Q _532_/Q VGND VGND VPWR VPWR _375_/B sky130_fd_sc_hd__xor2_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_354_ _523_/Q _526_/Q VGND VGND VPWR VPWR _358_/B sky130_fd_sc_hd__xor2_1
X_423_ _427_/A VGND VGND VPWR VPWR _423_/Y sky130_fd_sc_hd__inv_2
X_285_ _497_/Q _500_/Q VGND VGND VPWR VPWR _289_/B sky130_fd_sc_hd__xor2_1
Xinput7 x[14] VGND VGND VPWR VPWR _309_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_337_ _337_/A _337_/B VGND VGND VPWR VPWR _516_/D sky130_fd_sc_hd__xnor2_1
X_268_ _491_/Q _494_/Q VGND VGND VPWR VPWR _272_/B sky130_fd_sc_hd__xor2_1
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_406_ _409_/A VGND VGND VPWR VPWR _406_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput21 x[27] VGND VGND VPWR VPWR _379_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 x[17] VGND VGND VPWR VPWR _325_/B sky130_fd_sc_hd__clkbuf_1
Xinput32 x[8] VGND VGND VPWR VPWR _276_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_370_ _370_/A _370_/B VGND VGND VPWR VPWR _528_/D sky130_fd_sc_hd__xnor2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_499_ _505_/CLK _499_/D _427_/Y VGND VGND VPWR VPWR _499_/Q sky130_fd_sc_hd__dfrtp_1
X_353_ _353_/A _353_/B VGND VGND VPWR VPWR _522_/D sky130_fd_sc_hd__xnor2_1
X_284_ _394_/A VGND VGND VPWR VPWR _284_/X sky130_fd_sc_hd__clkbuf_2
X_422_ _428_/A VGND VGND VPWR VPWR _427_/A sky130_fd_sc_hd__buf_2
Xinput8 x[15] VGND VGND VPWR VPWR _315_/B sky130_fd_sc_hd__clkbuf_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_336_ _357_/A _336_/B VGND VGND VPWR VPWR _337_/A sky130_fd_sc_hd__nand2_1
X_267_ _267_/A _267_/B VGND VGND VPWR VPWR _490_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_405_ _409_/A VGND VGND VPWR VPWR _405_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput22 x[28] VGND VGND VPWR VPWR _384_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 x[18] VGND VGND VPWR VPWR _330_/B sky130_fd_sc_hd__clkbuf_1
Xinput33 x[9] VGND VGND VPWR VPWR _282_/B sky130_fd_sc_hd__clkbuf_1
X_319_ _311_/X _320_/B _321_/B _318_/X VGND VGND VPWR VPWR _509_/D sky130_fd_sc_hd__a31o_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_498_ _505_/CLK _498_/D _426_/Y VGND VGND VPWR VPWR _498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_421_ _421_/A VGND VGND VPWR VPWR _421_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 x[16] VGND VGND VPWR VPWR _320_/B sky130_fd_sc_hd__clkbuf_1
X_352_ _357_/A _352_/B VGND VGND VPWR VPWR _353_/A sky130_fd_sc_hd__nand2_1
X_283_ _283_/A _283_/B VGND VGND VPWR VPWR _496_/D sky130_fd_sc_hd__xnor2_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_266_ _276_/A _266_/B VGND VGND VPWR VPWR _267_/A sky130_fd_sc_hd__nand2_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_335_ _362_/A VGND VGND VPWR VPWR _357_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_404_ _428_/A VGND VGND VPWR VPWR _409_/A sky130_fd_sc_hd__buf_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput23 x[29] VGND VGND VPWR VPWR _389_/B sky130_fd_sc_hd__clkbuf_2
Xinput34 y VGND VGND VPWR VPWR _253_/A sky130_fd_sc_hd__clkbuf_2
Xinput12 x[19] VGND VGND VPWR VPWR _336_/B sky130_fd_sc_hd__clkbuf_1
X_318_ _509_/Q _512_/Q VGND VGND VPWR VPWR _318_/X sky130_fd_sc_hd__and2_1
X_249_ _249_/A _249_/B VGND VGND VPWR VPWR _484_/D sky130_fd_sc_hd__xnor2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_497_ _497_/CLK _497_/D _425_/Y VGND VGND VPWR VPWR _497_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_351_ _338_/X _352_/B _353_/B _350_/X VGND VGND VPWR VPWR _521_/D sky130_fd_sc_hd__a31o_1
X_420_ _421_/A VGND VGND VPWR VPWR _420_/Y sky130_fd_sc_hd__inv_2
X_282_ _303_/A _282_/B VGND VGND VPWR VPWR _283_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _311_/X _336_/B _337_/B _333_/X VGND VGND VPWR VPWR _515_/D sky130_fd_sc_hd__a31o_1
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_403_ _465_/A VGND VGND VPWR VPWR _428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_265_ _257_/X _266_/B _267_/B _264_/X VGND VGND VPWR VPWR _489_/D sky130_fd_sc_hd__a31o_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 x[2] VGND VGND VPWR VPWR _243_/B sky130_fd_sc_hd__clkbuf_2
Xinput13 x[1] VGND VGND VPWR VPWR _238_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_317_ _509_/Q _512_/Q VGND VGND VPWR VPWR _321_/B sky130_fd_sc_hd__xor2_1
X_248_ _248_/A _248_/B VGND VGND VPWR VPWR _249_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_496_ _512_/CLK _496_/D _424_/Y VGND VGND VPWR VPWR _496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ _521_/Q _524_/Q VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__and2_1
X_281_ _362_/A VGND VGND VPWR VPWR _303_/A sky130_fd_sc_hd__clkbuf_2
X_479_ _497_/CLK _479_/D _402_/Y VGND VGND VPWR VPWR _479_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ _489_/Q _492_/Q VGND VGND VPWR VPWR _264_/X sky130_fd_sc_hd__and2_1
X_333_ _515_/Q _518_/Q VGND VGND VPWR VPWR _333_/X sky130_fd_sc_hd__and2_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_402_ _402_/A VGND VGND VPWR VPWR _402_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput25 x[30] VGND VGND VPWR VPWR _394_/B sky130_fd_sc_hd__clkbuf_2
Xinput14 x[20] VGND VGND VPWR VPWR _342_/B sky130_fd_sc_hd__clkbuf_1
X_316_ _316_/A _316_/B VGND VGND VPWR VPWR _508_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_247_ _223_/X _248_/B _249_/B _246_/X VGND VGND VPWR VPWR _483_/D sky130_fd_sc_hd__a31o_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_495_ _497_/CLK _495_/D _423_/Y VGND VGND VPWR VPWR _495_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_280_ _257_/X _282_/B _283_/B _279_/X VGND VGND VPWR VPWR _495_/D sky130_fd_sc_hd__a31o_1
X_478_ _538_/CLK _478_/D _401_/Y VGND VGND VPWR VPWR _478_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ _489_/Q _492_/Q VGND VGND VPWR VPWR _267_/B sky130_fd_sc_hd__xor2_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _515_/Q _518_/Q VGND VGND VPWR VPWR _337_/B sky130_fd_sc_hd__xor2_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_401_ _402_/A VGND VGND VPWR VPWR _401_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 x[31] VGND VGND VPWR VPWR _232_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 x[21] VGND VGND VPWR VPWR _347_/B sky130_fd_sc_hd__clkbuf_1
X_315_ _330_/A _315_/B VGND VGND VPWR VPWR _316_/A sky130_fd_sc_hd__nand2_1
X_246_ _483_/Q _486_/Q VGND VGND VPWR VPWR _246_/X sky130_fd_sc_hd__and2_1
XFILLER_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_229_ _248_/A _229_/B VGND VGND VPWR VPWR _230_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_494_ _512_/CLK _494_/D _421_/Y VGND VGND VPWR VPWR _494_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_477_ _536_/CLK _477_/D _400_/Y VGND VGND VPWR VPWR _477_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _331_/A _331_/B VGND VGND VPWR VPWR _514_/D sky130_fd_sc_hd__xnor2_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_262_ _262_/A _262_/B VGND VGND VPWR VPWR _488_/D sky130_fd_sc_hd__xnor2_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_400_ _402_/A VGND VGND VPWR VPWR _400_/Y sky130_fd_sc_hd__inv_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_529_ _536_/CLK _529_/D _464_/Y VGND VGND VPWR VPWR _529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput27 x[3] VGND VGND VPWR VPWR _248_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput16 x[22] VGND VGND VPWR VPWR _352_/B sky130_fd_sc_hd__clkbuf_1
X_314_ _311_/X _315_/B _316_/B _313_/X VGND VGND VPWR VPWR _507_/D sky130_fd_sc_hd__a31o_1
X_245_ _483_/Q _486_/Q VGND VGND VPWR VPWR _249_/B sky130_fd_sc_hd__xor2_1
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_228_ _365_/A VGND VGND VPWR VPWR _248_/A sky130_fd_sc_hd__buf_2
XFILLER_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_493_ _493_/CLK _493_/D _420_/Y VGND VGND VPWR VPWR _493_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_476_ _497_/CLK _476_/D _399_/Y VGND VGND VPWR VPWR _476_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _330_/A _330_/B VGND VGND VPWR VPWR _331_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _276_/A _261_/B VGND VGND VPWR VPWR _262_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_459_ _459_/A VGND VGND VPWR VPWR _464_/A sky130_fd_sc_hd__buf_2
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_528_ _536_/CLK _528_/D _463_/Y VGND VGND VPWR VPWR _528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 x[4] VGND VGND VPWR VPWR _255_/B sky130_fd_sc_hd__clkbuf_1
Xinput17 x[23] VGND VGND VPWR VPWR _357_/B sky130_fd_sc_hd__clkbuf_1
X_313_ _507_/Q _510_/Q VGND VGND VPWR VPWR _313_/X sky130_fd_sc_hd__and2_1
X_244_ _244_/A _244_/B VGND VGND VPWR VPWR _482_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ _253_/A VGND VGND VPWR VPWR _365_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_492_ _512_/CLK _492_/D _419_/Y VGND VGND VPWR VPWR _492_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_475_ _497_/CLK _475_/D _398_/Y VGND VGND VPWR VPWR _475_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_260_ _257_/X _261_/B _262_/B _259_/X VGND VGND VPWR VPWR _487_/D sky130_fd_sc_hd__a31o_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_458_ _458_/A VGND VGND VPWR VPWR _458_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_527_ _536_/CLK _527_/D _462_/Y VGND VGND VPWR VPWR _527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_389_ _394_/A _389_/B VGND VGND VPWR VPWR _390_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput29 x[5] VGND VGND VPWR VPWR _261_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 x[24] VGND VGND VPWR VPWR _363_/B sky130_fd_sc_hd__clkbuf_1
X_312_ _507_/Q _510_/Q VGND VGND VPWR VPWR _316_/B sky130_fd_sc_hd__xor2_1
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_243_ _248_/A _243_/B VGND VGND VPWR VPWR _244_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_226_ _223_/X _229_/B _230_/B _225_/X VGND VGND VPWR VPWR _475_/D sky130_fd_sc_hd__a31o_1
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_491_ _512_/CLK _491_/D _418_/Y VGND VGND VPWR VPWR _491_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_474_ _474_/A VGND VGND VPWR VPWR _474_/Y sky130_fd_sc_hd__inv_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_526_ _526_/CLK _526_/D _461_/Y VGND VGND VPWR VPWR _526_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_457_ _458_/A VGND VGND VPWR VPWR _457_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_388_ _365_/X _389_/B _390_/B _387_/X VGND VGND VPWR VPWR _535_/D sky130_fd_sc_hd__a31o_1
Xinput19 x[25] VGND VGND VPWR VPWR _369_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_311_ _365_/A VGND VGND VPWR VPWR _311_/X sky130_fd_sc_hd__clkbuf_2
X_242_ _223_/X _243_/B _244_/B _241_/X VGND VGND VPWR VPWR _481_/D sky130_fd_sc_hd__a31o_1
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_509_ _518_/CLK _509_/D _440_/Y VGND VGND VPWR VPWR _509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_225_ _475_/Q _480_/Q VGND VGND VPWR VPWR _225_/X sky130_fd_sc_hd__and2_1
XFILLER_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_490_ _493_/CLK _490_/D _417_/Y VGND VGND VPWR VPWR _490_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_473_ _474_/A VGND VGND VPWR VPWR _473_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR _526_/CLK sky130_fd_sc_hd__clkbuf_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_456_ _458_/A VGND VGND VPWR VPWR _456_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_525_ _536_/CLK _525_/D _460_/Y VGND VGND VPWR VPWR _525_/Q sky130_fd_sc_hd__dfrtp_1
X_387_ _535_/Q _538_/Q VGND VGND VPWR VPWR _387_/X sky130_fd_sc_hd__and2_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_310_ _310_/A _310_/B VGND VGND VPWR VPWR _506_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_439_ _440_/A VGND VGND VPWR VPWR _439_/Y sky130_fd_sc_hd__inv_2
X_508_ _538_/CLK _508_/D _439_/Y VGND VGND VPWR VPWR _508_/Q sky130_fd_sc_hd__dfrtp_1
X_241_ _481_/Q _484_/Q VGND VGND VPWR VPWR _241_/X sky130_fd_sc_hd__and2_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_224_ _475_/Q _480_/Q VGND VGND VPWR VPWR _230_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_472_ _474_/A VGND VGND VPWR VPWR _472_/Y sky130_fd_sc_hd__inv_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_455_ _458_/A VGND VGND VPWR VPWR _455_/Y sky130_fd_sc_hd__inv_2
X_524_ _526_/CLK _524_/D _458_/Y VGND VGND VPWR VPWR _524_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_386_ _535_/Q _538_/Q VGND VGND VPWR VPWR _390_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR _518_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_240_ _481_/Q _484_/Q VGND VGND VPWR VPWR _244_/B sky130_fd_sc_hd__xor2_1
X_507_ _518_/CLK _507_/D _438_/Y VGND VGND VPWR VPWR _507_/Q sky130_fd_sc_hd__dfrtp_1
X_438_ _440_/A VGND VGND VPWR VPWR _438_/Y sky130_fd_sc_hd__inv_2
X_369_ _384_/A _369_/B VGND VGND VPWR VPWR _370_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_223_ _394_/A VGND VGND VPWR VPWR _223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_471_ _474_/A VGND VGND VPWR VPWR _471_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_454_ _458_/A VGND VGND VPWR VPWR _454_/Y sky130_fd_sc_hd__inv_2
X_523_ _526_/CLK _523_/D _457_/Y VGND VGND VPWR VPWR _523_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_385_ _385_/A _385_/B VGND VGND VPWR VPWR _534_/D sky130_fd_sc_hd__xnor2_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_368_ _365_/X _369_/B _370_/B _367_/X VGND VGND VPWR VPWR _527_/D sky130_fd_sc_hd__a31o_1
X_437_ _440_/A VGND VGND VPWR VPWR _437_/Y sky130_fd_sc_hd__inv_2
X_299_ _299_/A _299_/B VGND VGND VPWR VPWR _502_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_506_ _538_/CLK _506_/D _437_/Y VGND VGND VPWR VPWR _506_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_222_ _253_/A VGND VGND VPWR VPWR _394_/A sky130_fd_sc_hd__buf_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR _536_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_470_ _470_/A VGND VGND VPWR VPWR _470_/Y sky130_fd_sc_hd__inv_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_522_ _526_/CLK _522_/D _456_/Y VGND VGND VPWR VPWR _522_/Q sky130_fd_sc_hd__dfrtp_1
X_453_ _459_/A VGND VGND VPWR VPWR _458_/A sky130_fd_sc_hd__buf_2
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_384_ _384_/A _384_/B VGND VGND VPWR VPWR _385_/A sky130_fd_sc_hd__nand2_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_367_ _527_/Q _530_/Q VGND VGND VPWR VPWR _367_/X sky130_fd_sc_hd__and2_1
X_505_ _505_/CLK _505_/D _436_/Y VGND VGND VPWR VPWR _505_/Q sky130_fd_sc_hd__dfrtp_1
X_436_ _440_/A VGND VGND VPWR VPWR _436_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ _303_/A _298_/B VGND VGND VPWR VPWR _299_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_419_ _421_/A VGND VGND VPWR VPWR _419_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR _538_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_521_ _526_/CLK _521_/D _455_/Y VGND VGND VPWR VPWR _521_/Q sky130_fd_sc_hd__dfrtp_1
X_452_ _452_/A VGND VGND VPWR VPWR _452_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _365_/X _384_/B _385_/B _382_/X VGND VGND VPWR VPWR _533_/D sky130_fd_sc_hd__a31o_1
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_366_ _527_/Q _530_/Q VGND VGND VPWR VPWR _370_/B sky130_fd_sc_hd__xor2_1
X_435_ _459_/A VGND VGND VPWR VPWR _440_/A sky130_fd_sc_hd__buf_2
X_504_ _538_/CLK _504_/D _433_/Y VGND VGND VPWR VPWR _504_/Q sky130_fd_sc_hd__dfrtp_1
X_297_ _284_/X _298_/B _299_/B _296_/X VGND VGND VPWR VPWR _501_/D sky130_fd_sc_hd__a31o_1
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_418_ _421_/A VGND VGND VPWR VPWR _418_/Y sky130_fd_sc_hd__inv_2
X_349_ _521_/Q _524_/Q VGND VGND VPWR VPWR _353_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_520_ _526_/CLK _520_/D _454_/Y VGND VGND VPWR VPWR _520_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_451_ _452_/A VGND VGND VPWR VPWR _451_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR _512_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_382_ _533_/Q _536_/Q VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__and2_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_365_ _365_/A VGND VGND VPWR VPWR _365_/X sky130_fd_sc_hd__clkbuf_2
X_434_ _465_/A VGND VGND VPWR VPWR _459_/A sky130_fd_sc_hd__clkbuf_2
X_296_ _501_/Q _504_/Q VGND VGND VPWR VPWR _296_/X sky130_fd_sc_hd__and2_1
X_503_ _505_/CLK _503_/D _432_/Y VGND VGND VPWR VPWR _503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_417_ _421_/A VGND VGND VPWR VPWR _417_/Y sky130_fd_sc_hd__inv_2
X_348_ _348_/A _348_/B VGND VGND VPWR VPWR _520_/D sky130_fd_sc_hd__xnor2_1
X_279_ _495_/Q _498_/Q VGND VGND VPWR VPWR _279_/X sky130_fd_sc_hd__and2_1
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_450_ _452_/A VGND VGND VPWR VPWR _450_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_381_ _533_/Q _536_/Q VGND VGND VPWR VPWR _385_/B sky130_fd_sc_hd__xor2_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_433_ _433_/A VGND VGND VPWR VPWR _433_/Y sky130_fd_sc_hd__inv_2
X_502_ _505_/CLK _502_/D _431_/Y VGND VGND VPWR VPWR _502_/Q sky130_fd_sc_hd__dfrtp_1
X_364_ _364_/A _364_/B VGND VGND VPWR VPWR _526_/D sky130_fd_sc_hd__xnor2_1
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_295_ _501_/Q _504_/Q VGND VGND VPWR VPWR _299_/B sky130_fd_sc_hd__xor2_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR _493_/CLK sky130_fd_sc_hd__clkbuf_2
X_347_ _357_/A _347_/B VGND VGND VPWR VPWR _348_/A sky130_fd_sc_hd__nand2_1
X_416_ _428_/A VGND VGND VPWR VPWR _421_/A sky130_fd_sc_hd__buf_2
X_278_ _495_/Q _498_/Q VGND VGND VPWR VPWR _283_/B sky130_fd_sc_hd__xor2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_380_ _380_/A _380_/B VGND VGND VPWR VPWR _532_/D sky130_fd_sc_hd__xnor2_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

